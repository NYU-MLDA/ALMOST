//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n986_, new_n987_,
    new_n989_, new_n990_, new_n991_, new_n993_, new_n994_, new_n995_,
    new_n997_, new_n998_, new_n999_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1028_, new_n1029_, new_n1031_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1046_,
    new_n1047_, new_n1048_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1055_, new_n1056_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT6), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(KEYINPUT9), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n205_), .A2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G85gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n211_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n208_), .A2(new_n209_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n204_), .B(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n213_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n220_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n221_), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n226_), .B(new_n225_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n220_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n219_), .B1(new_n229_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G64gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G78gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(KEYINPUT11), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G78gat), .Z(new_n239_));
  INV_X1    g038(.A(G64gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G57gat), .ZN(new_n241_));
  INV_X1    g040(.A(G57gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G64gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n243_), .A3(KEYINPUT11), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n238_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n203_), .B1(new_n235_), .B2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n211_), .A2(new_n218_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n234_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n233_), .B1(new_n232_), .B2(new_n220_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n247_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT66), .A3(new_n253_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n249_), .B(new_n247_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n235_), .A2(KEYINPUT65), .A3(new_n247_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n248_), .A2(new_n254_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(new_n235_), .B2(new_n247_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n261_), .B1(new_n235_), .B2(new_n247_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n252_), .A2(new_n253_), .A3(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G120gat), .B(G148gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT5), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G176gat), .B(G204gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n270_), .B(new_n271_), .Z(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n262_), .A2(new_n268_), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n262_), .B2(new_n268_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n262_), .A2(new_n268_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n272_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n262_), .A2(new_n268_), .A3(new_n273_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT68), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n202_), .B1(new_n277_), .B2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n276_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(KEYINPUT68), .A3(new_n280_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT13), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n282_), .A2(KEYINPUT69), .A3(new_n285_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G113gat), .B(G141gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT77), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G169gat), .B(G197gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G43gat), .B(G50gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G29gat), .B(G36gat), .Z(new_n300_));
  XOR2_X1   g099(.A(G43gat), .B(G50gat), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G15gat), .B(G22gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G1gat), .A2(G8gat), .ZN(new_n304_));
  INV_X1    g103(.A(G1gat), .ZN(new_n305_));
  INV_X1    g104(.A(G8gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(KEYINPUT14), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n303_), .A2(new_n304_), .A3(new_n307_), .A4(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n303_), .A2(new_n308_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n299_), .B(new_n302_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(new_n299_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n311_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n309_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n315_), .A3(KEYINPUT76), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G229gat), .A2(G233gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n309_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n299_), .A4(new_n302_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n316_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT15), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n313_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n302_), .A2(KEYINPUT15), .A3(new_n299_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n319_), .A3(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n317_), .A3(new_n315_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n296_), .B1(new_n322_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n327_), .A3(new_n296_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(KEYINPUT78), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n330_), .B2(KEYINPUT78), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n329_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(KEYINPUT78), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT79), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT25), .B(G183gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT80), .B1(new_n341_), .B2(G190gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G190gat), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n340_), .B(new_n342_), .C1(new_n343_), .C2(KEYINPUT80), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT24), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT81), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n352_), .A2(G169gat), .A3(G176gat), .ZN(new_n353_));
  INV_X1    g152(.A(G169gat), .ZN(new_n354_));
  INV_X1    g153(.A(G176gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT81), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n351_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n355_), .A3(KEYINPUT81), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n352_), .B1(G169gat), .B2(G176gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(KEYINPUT24), .A4(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n344_), .A2(new_n350_), .A3(new_n357_), .A4(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G183gat), .ZN(new_n363_));
  INV_X1    g162(.A(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n347_), .A2(new_n348_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n360_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT82), .B(G176gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT22), .B(G169gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n366_), .B1(new_n370_), .B2(KEYINPUT83), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n372_));
  AOI211_X1 g171(.A(new_n372_), .B(new_n367_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n362_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT30), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G71gat), .B(G99gat), .ZN(new_n377_));
  INV_X1    g176(.A(G43gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(G15gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n379_), .B(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n375_), .A2(new_n376_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n375_), .A2(new_n376_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n383_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n375_), .A2(new_n376_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n384_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT86), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n384_), .B(new_n391_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G113gat), .B(G120gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G134gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G127gat), .ZN(new_n396_));
  INV_X1    g195(.A(G127gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G134gat), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n396_), .A2(new_n398_), .A3(KEYINPUT85), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT85), .B1(new_n396_), .B2(new_n398_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n394_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n398_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n396_), .A2(new_n398_), .A3(KEYINPUT85), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n393_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT31), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n390_), .A2(new_n392_), .A3(new_n408_), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n389_), .A2(KEYINPUT86), .A3(new_n408_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT99), .ZN(new_n412_));
  XOR2_X1   g211(.A(G8gat), .B(G36gat), .Z(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT18), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G226gat), .A2(G233gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT19), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n355_), .A2(KEYINPUT82), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G176gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n354_), .A2(KEYINPUT22), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT22), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G169gat), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n360_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n428_), .A2(new_n372_), .B1(new_n350_), .B2(new_n365_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n373_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n363_), .A2(KEYINPUT25), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT25), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G183gat), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n342_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n364_), .A2(KEYINPUT26), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n341_), .A2(G190gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n353_), .A2(new_n356_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n367_), .A2(new_n351_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n434_), .A2(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT24), .B1(new_n358_), .B2(new_n359_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(new_n349_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n429_), .A2(new_n430_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT91), .ZN(new_n446_));
  INV_X1    g245(.A(G197gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(G204gat), .ZN(new_n448_));
  INV_X1    g247(.A(G204gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(G204gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT21), .ZN(new_n453_));
  INV_X1    g252(.A(G218gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G211gat), .ZN(new_n455_));
  INV_X1    g254(.A(G211gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G218gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n453_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n452_), .A2(new_n458_), .A3(KEYINPUT92), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n455_), .A2(new_n457_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n449_), .A2(G197gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n451_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(KEYINPUT21), .B2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n448_), .A2(new_n450_), .A3(new_n453_), .A4(new_n451_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n461_), .A2(new_n462_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT95), .B1(new_n445_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n467_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n462_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT92), .B1(new_n452_), .B2(new_n458_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT95), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n374_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n366_), .A2(KEYINPUT94), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n347_), .A2(new_n365_), .A3(new_n479_), .A4(new_n348_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n428_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n435_), .A2(new_n436_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n361_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n357_), .A2(new_n350_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(KEYINPUT93), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT93), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n357_), .A2(new_n486_), .A3(new_n350_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n481_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n477_), .B1(new_n488_), .B2(new_n468_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n420_), .B1(new_n476_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT20), .B1(new_n374_), .B2(new_n473_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT93), .B1(new_n443_), .B2(new_n349_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n487_), .A2(new_n492_), .A3(new_n482_), .A4(new_n361_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n478_), .A2(new_n480_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n370_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n461_), .A2(new_n462_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n493_), .A2(new_n495_), .B1(new_n496_), .B2(new_n470_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n491_), .A2(new_n497_), .A3(new_n419_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n412_), .B(new_n417_), .C1(new_n490_), .C2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n468_), .A2(new_n495_), .A3(new_n493_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n419_), .A2(new_n477_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n493_), .A2(new_n495_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n473_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n429_), .A2(new_n430_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(new_n468_), .A3(new_n362_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(KEYINPUT20), .A3(new_n507_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n476_), .A2(new_n503_), .B1(new_n508_), .B2(new_n419_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT99), .B1(new_n509_), .B2(new_n416_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n475_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n474_), .B1(new_n374_), .B2(new_n473_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n489_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n419_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n498_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n416_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(KEYINPUT27), .B(new_n499_), .C1(new_n510_), .C2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT29), .ZN(new_n518_));
  OR2_X1    g317(.A1(G141gat), .A2(G148gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G141gat), .A2(G148gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G155gat), .A2(G162gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G155gat), .A2(G162gat), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(KEYINPUT1), .B2(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(KEYINPUT1), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n521_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT3), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT3), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT87), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G141gat), .A2(G148gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n520_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT2), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT2), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n520_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n532_), .A2(new_n535_), .A3(new_n536_), .A4(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n540_));
  AND2_X1   g339(.A1(G155gat), .A2(G162gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n540_), .B1(new_n541_), .B2(new_n522_), .ZN(new_n542_));
  INV_X1    g341(.A(G155gat), .ZN(new_n543_));
  INV_X1    g342(.A(G162gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(KEYINPUT89), .A3(new_n523_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n526_), .B1(new_n539_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n473_), .B1(new_n518_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G106gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n539_), .A2(new_n547_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n526_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G22gat), .B(G50gat), .ZN(new_n555_));
  AND4_X1   g354(.A1(new_n518_), .A2(new_n553_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n548_), .B2(new_n518_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n552_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n553_), .A2(new_n518_), .A3(new_n554_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n555_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n548_), .A2(new_n518_), .A3(new_n555_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n551_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G228gat), .A2(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(G78gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n558_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n558_), .B2(new_n563_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n550_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n556_), .A2(new_n557_), .A3(new_n552_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n551_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n566_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n549_), .B(new_n213_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n558_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT27), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n502_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n477_), .B1(new_n445_), .B2(new_n468_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n420_), .B1(new_n581_), .B2(new_n505_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n580_), .A2(new_n582_), .A3(new_n417_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n500_), .B(new_n501_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n419_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n416_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n579_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n517_), .A2(new_n578_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n553_), .A2(new_n554_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n401_), .A2(new_n406_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n548_), .A2(new_n407_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G225gat), .A2(G233gat), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n591_), .A2(KEYINPUT4), .A3(new_n592_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n593_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n591_), .B2(KEYINPUT4), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n594_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G1gat), .B(G29gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G57gat), .B(G85gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n594_), .B(new_n605_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n411_), .A2(new_n588_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n592_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n548_), .A2(new_n407_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT4), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n593_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n591_), .A2(KEYINPUT4), .A3(new_n592_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n613_), .A2(new_n593_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n603_), .A2(new_n609_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT97), .B1(new_n611_), .B2(new_n612_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n591_), .A2(new_n621_), .A3(new_n592_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n596_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n596_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n605_), .B1(new_n624_), .B2(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n610_), .A2(new_n619_), .A3(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n583_), .A2(new_n586_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n610_), .A2(new_n619_), .A3(new_n626_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n417_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n584_), .A2(new_n585_), .A3(new_n416_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT98), .B1(new_n631_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n416_), .A2(KEYINPUT32), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n509_), .A2(new_n636_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n500_), .A2(KEYINPUT20), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n515_), .B1(new_n639_), .B2(new_n420_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(KEYINPUT32), .A3(new_n416_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n630_), .A2(new_n635_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n578_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n640_), .A2(new_n417_), .B1(new_n633_), .B2(new_n412_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n498_), .B1(new_n513_), .B2(new_n419_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(KEYINPUT99), .A3(new_n416_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n646_), .A2(new_n648_), .A3(new_n579_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n607_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n577_), .A2(new_n587_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n645_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n570_), .A2(new_n576_), .A3(new_n604_), .A4(new_n606_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT27), .B1(new_n632_), .B2(new_n633_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(KEYINPUT100), .A3(new_n517_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n644_), .A2(new_n652_), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n608_), .B1(new_n657_), .B2(new_n411_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n291_), .A2(new_n339_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(G231gat), .A2(G233gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n247_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT72), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n241_), .A2(new_n243_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT11), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n244_), .A3(new_n239_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n660_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n238_), .A3(new_n667_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n661_), .A2(new_n662_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n662_), .B1(new_n661_), .B2(new_n668_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n319_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n668_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n667_), .B1(new_n666_), .B2(new_n238_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT72), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n319_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n661_), .A2(new_n662_), .A3(new_n668_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(G127gat), .B(G155gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(G183gat), .B(G211gat), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n678_), .B(new_n679_), .Z(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n682_), .A2(new_n683_), .A3(KEYINPUT17), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT17), .B1(new_n682_), .B2(new_n683_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n671_), .A2(new_n677_), .A3(new_n684_), .A4(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n671_), .B2(new_n677_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT74), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT74), .B(new_n685_), .C1(new_n671_), .C2(new_n677_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT75), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n686_), .B(KEYINPUT75), .C1(new_n689_), .C2(new_n690_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT37), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n252_), .A2(new_n325_), .A3(new_n324_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n235_), .A2(new_n313_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n700_));
  NAND2_X1  g499(.A1(G232gat), .A2(G233gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT35), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n699_), .A3(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n702_), .A2(new_n703_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(G190gat), .B(G218gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(G134gat), .B(G162gat), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(KEYINPUT36), .ZN(new_n711_));
  INV_X1    g510(.A(new_n706_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n698_), .A2(new_n699_), .A3(new_n712_), .A4(new_n704_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n707_), .A2(new_n711_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n710_), .B(KEYINPUT36), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n707_), .B2(new_n713_), .ZN(new_n717_));
  OAI211_X1 g516(.A(KEYINPUT71), .B(new_n697_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n707_), .A2(new_n713_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n697_), .A2(KEYINPUT71), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n697_), .A2(KEYINPUT71), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n721_), .A2(new_n714_), .A3(new_n722_), .A4(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n718_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n696_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n659_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT101), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n659_), .A2(new_n730_), .A3(new_n727_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n305_), .A3(new_n607_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT38), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n732_), .A2(KEYINPUT38), .A3(new_n305_), .A4(new_n607_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n339_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n288_), .A2(new_n695_), .A3(new_n289_), .A4(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n715_), .A2(new_n717_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n738_), .A2(new_n658_), .A3(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G1gat), .B1(new_n741_), .B2(new_n650_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n735_), .A2(new_n736_), .A3(new_n742_), .ZN(G1324gat));
  NAND2_X1  g542(.A1(new_n517_), .A2(new_n587_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n729_), .A2(new_n306_), .A3(new_n744_), .A4(new_n731_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n744_), .ZN(new_n746_));
  NOR4_X1   g545(.A1(new_n738_), .A2(new_n658_), .A3(new_n739_), .A4(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n306_), .B1(new_n747_), .B2(KEYINPUT102), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n740_), .A2(new_n744_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n748_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n748_), .B2(new_n751_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n745_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT40), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI211_X1 g556(.A(KEYINPUT40), .B(new_n745_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1325gat));
  INV_X1    g558(.A(new_n411_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n740_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G15gat), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT104), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT104), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT41), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n732_), .A2(new_n381_), .A3(new_n760_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n763_), .A2(KEYINPUT41), .A3(new_n764_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(G1326gat));
  INV_X1    g569(.A(G22gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n732_), .A2(new_n771_), .A3(new_n577_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n740_), .B2(new_n577_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT42), .Z(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1327gat));
  INV_X1    g574(.A(new_n739_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n695_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n659_), .A2(new_n777_), .ZN(new_n778_));
  OR3_X1    g577(.A1(new_n778_), .A2(G29gat), .A3(new_n650_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n290_), .A2(new_n696_), .A3(new_n737_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n781_));
  INV_X1    g580(.A(new_n608_), .ZN(new_n782_));
  AOI22_X1  g581(.A1(new_n617_), .A2(new_n618_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n783_), .A2(new_n633_), .A3(new_n632_), .A4(new_n610_), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n784_), .A2(KEYINPUT98), .B1(new_n637_), .B2(new_n641_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n577_), .B1(new_n785_), .B2(new_n630_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n655_), .A2(KEYINPUT100), .A3(new_n517_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT100), .B1(new_n655_), .B2(new_n517_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n782_), .B1(new_n789_), .B2(new_n760_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n781_), .B1(new_n790_), .B2(new_n726_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n658_), .A2(KEYINPUT43), .A3(new_n725_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT44), .B(new_n780_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n290_), .A2(new_n696_), .A3(new_n737_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT43), .B1(new_n658_), .B2(new_n725_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n655_), .A2(new_n517_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n578_), .A2(new_n643_), .B1(new_n798_), .B2(new_n645_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n760_), .B1(new_n799_), .B2(new_n656_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n781_), .B(new_n726_), .C1(new_n800_), .C2(new_n608_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n796_), .B1(new_n797_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n795_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n805_));
  INV_X1    g604(.A(new_n802_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n650_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(new_n805_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(G29gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n805_), .B1(new_n804_), .B2(new_n809_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n779_), .B1(new_n811_), .B2(new_n812_), .ZN(G1328gat));
  INV_X1    g612(.A(KEYINPUT46), .ZN(new_n814_));
  INV_X1    g613(.A(G36gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n744_), .B1(new_n802_), .B2(new_n807_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n804_), .B2(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n659_), .A2(new_n777_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n744_), .B(KEYINPUT108), .Z(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(G36gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n822_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT45), .B1(new_n778_), .B2(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n814_), .B1(new_n818_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n825_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n816_), .B1(new_n795_), .B2(new_n803_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT46), .B(new_n828_), .C1(new_n829_), .C2(new_n815_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(G1329gat));
  NAND2_X1  g630(.A1(new_n806_), .A2(new_n808_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n411_), .A2(new_n378_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n793_), .A2(new_n794_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT106), .B1(new_n802_), .B2(KEYINPUT44), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n832_), .B(new_n833_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n378_), .B1(new_n778_), .B2(new_n411_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n836_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1330gat));
  AOI21_X1  g642(.A(G50gat), .B1(new_n819_), .B2(new_n577_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n804_), .A2(new_n832_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n577_), .A2(G50gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(G1331gat));
  NAND3_X1  g646(.A1(new_n693_), .A2(new_n339_), .A3(new_n694_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n290_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n658_), .A2(new_n739_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G57gat), .B1(new_n851_), .B2(new_n650_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n790_), .A2(new_n339_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n853_), .A2(KEYINPUT110), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n290_), .B1(new_n853_), .B2(KEYINPUT110), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n727_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n607_), .A2(new_n242_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n852_), .B1(new_n856_), .B2(new_n857_), .ZN(G1332gat));
  OAI21_X1  g657(.A(G64gat), .B1(new_n851_), .B2(new_n821_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT48), .ZN(new_n860_));
  INV_X1    g659(.A(new_n821_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n240_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n856_), .B2(new_n862_), .ZN(G1333gat));
  OAI21_X1  g662(.A(G71gat), .B1(new_n851_), .B2(new_n411_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n866_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n411_), .A2(G71gat), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n867_), .A2(new_n868_), .B1(new_n856_), .B2(new_n869_), .ZN(G1334gat));
  NAND2_X1  g669(.A1(new_n577_), .A2(new_n565_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n856_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G78gat), .B1(new_n851_), .B2(new_n578_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(KEYINPUT50), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(KEYINPUT50), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n872_), .B(KEYINPUT112), .C1(new_n874_), .C2(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1335gat));
  NAND2_X1  g679(.A1(new_n797_), .A2(new_n801_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n290_), .A2(new_n695_), .A3(new_n737_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n883_), .A2(new_n216_), .A3(new_n650_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n854_), .A2(new_n777_), .A3(new_n855_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n206_), .B1(new_n885_), .B2(new_n650_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n887_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n884_), .B1(new_n888_), .B2(new_n889_), .ZN(G1336gat));
  OAI21_X1  g689(.A(G92gat), .B1(new_n883_), .B2(new_n821_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n744_), .A2(new_n207_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n885_), .B2(new_n892_), .ZN(G1337gat));
  NAND2_X1  g692(.A1(new_n212_), .A2(new_n214_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n885_), .A2(new_n894_), .A3(new_n411_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n883_), .A2(new_n411_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n224_), .ZN(new_n897_));
  OR3_X1    g696(.A1(new_n895_), .A2(new_n897_), .A3(KEYINPUT51), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT51), .B1(new_n895_), .B2(new_n897_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1338gat));
  NAND3_X1  g699(.A1(new_n881_), .A2(new_n577_), .A3(new_n882_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n901_), .A2(G106gat), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n901_), .B2(G106gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n577_), .A2(new_n213_), .ZN(new_n905_));
  OAI22_X1  g704(.A1(new_n903_), .A2(new_n904_), .B1(new_n885_), .B2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT53), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n908_));
  OAI221_X1 g707(.A(new_n908_), .B1(new_n885_), .B2(new_n905_), .C1(new_n903_), .C2(new_n904_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1339gat));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n316_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n326_), .A2(new_n318_), .A3(new_n315_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(new_n295_), .A3(new_n913_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n914_), .A2(new_n330_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n283_), .A2(new_n284_), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n335_), .A2(new_n338_), .A3(new_n280_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT55), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n268_), .A2(new_n919_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .A4(KEYINPUT55), .ZN(new_n921_));
  AND4_X1   g720(.A1(new_n257_), .A2(new_n264_), .A3(new_n267_), .A4(new_n258_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n920_), .B(new_n921_), .C1(new_n922_), .C2(new_n260_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n272_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n923_), .A2(KEYINPUT56), .A3(new_n272_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n918_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n776_), .B1(new_n917_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT57), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n280_), .A2(new_n915_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n725_), .B1(new_n932_), .B2(KEYINPUT58), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n926_), .A2(new_n927_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n929_), .A2(new_n930_), .B1(new_n933_), .B2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n934_), .A2(new_n280_), .A3(new_n737_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n739_), .B1(new_n940_), .B2(new_n916_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(KEYINPUT57), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n695_), .B1(new_n939_), .B2(new_n942_), .ZN(new_n943_));
  AND3_X1   g742(.A1(new_n693_), .A2(new_n694_), .A3(new_n339_), .ZN(new_n944_));
  AOI21_X1  g743(.A(KEYINPUT115), .B1(new_n286_), .B2(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT115), .ZN(new_n946_));
  AOI211_X1 g745(.A(new_n946_), .B(new_n848_), .C1(new_n282_), .C2(new_n285_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n725_), .B1(new_n945_), .B2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(KEYINPUT54), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT13), .ZN(new_n950_));
  AOI21_X1  g749(.A(KEYINPUT13), .B1(new_n283_), .B2(new_n284_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n944_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n946_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n286_), .A2(KEYINPUT115), .A3(new_n944_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n955_), .A2(new_n956_), .A3(new_n725_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n943_), .B1(new_n949_), .B2(new_n957_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n411_), .A2(new_n588_), .A3(new_n650_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n911_), .B1(new_n958_), .B2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n933_), .A2(new_n938_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n962_), .B1(new_n941_), .B2(KEYINPUT57), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n929_), .A2(new_n930_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n696_), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n956_), .B1(new_n955_), .B2(new_n725_), .ZN(new_n966_));
  AOI211_X1 g765(.A(KEYINPUT54), .B(new_n726_), .C1(new_n953_), .C2(new_n954_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n968_), .A2(KEYINPUT59), .A3(new_n959_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n961_), .A2(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  OAI21_X1  g770(.A(G113gat), .B1(new_n971_), .B2(new_n339_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n958_), .A2(new_n960_), .ZN(new_n973_));
  INV_X1    g772(.A(G113gat), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n973_), .A2(new_n974_), .A3(new_n737_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n972_), .A2(new_n975_), .ZN(G1340gat));
  INV_X1    g775(.A(G120gat), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n977_), .B1(new_n290_), .B2(KEYINPUT60), .ZN(new_n978_));
  OAI211_X1 g777(.A(new_n973_), .B(new_n978_), .C1(KEYINPUT60), .C2(new_n977_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n290_), .B1(new_n961_), .B2(new_n969_), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n979_), .B1(new_n980_), .B2(new_n977_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n981_), .A2(KEYINPUT116), .ZN(new_n982_));
  INV_X1    g781(.A(KEYINPUT116), .ZN(new_n983_));
  OAI211_X1 g782(.A(new_n983_), .B(new_n979_), .C1(new_n980_), .C2(new_n977_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n982_), .A2(new_n984_), .ZN(G1341gat));
  OAI21_X1  g784(.A(G127gat), .B1(new_n971_), .B2(new_n696_), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n973_), .A2(new_n397_), .A3(new_n695_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n986_), .A2(new_n987_), .ZN(G1342gat));
  AOI21_X1  g787(.A(G134gat), .B1(new_n973_), .B2(new_n739_), .ZN(new_n989_));
  NOR2_X1   g788(.A1(new_n725_), .A2(new_n395_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n990_), .B(KEYINPUT117), .ZN(new_n991_));
  AOI21_X1  g790(.A(new_n989_), .B1(new_n970_), .B2(new_n991_), .ZN(G1343gat));
  NOR2_X1   g791(.A1(new_n958_), .A2(new_n760_), .ZN(new_n993_));
  NOR3_X1   g792(.A1(new_n861_), .A2(new_n578_), .A3(new_n650_), .ZN(new_n994_));
  NAND3_X1  g793(.A1(new_n993_), .A2(new_n737_), .A3(new_n994_), .ZN(new_n995_));
  XNOR2_X1  g794(.A(new_n995_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g795(.A1(new_n993_), .A2(new_n994_), .ZN(new_n997_));
  NOR2_X1   g796(.A1(new_n997_), .A2(new_n290_), .ZN(new_n998_));
  XOR2_X1   g797(.A(KEYINPUT118), .B(G148gat), .Z(new_n999_));
  XNOR2_X1  g798(.A(new_n998_), .B(new_n999_), .ZN(G1345gat));
  NAND4_X1  g799(.A1(new_n968_), .A2(new_n695_), .A3(new_n411_), .A4(new_n994_), .ZN(new_n1001_));
  OR2_X1    g800(.A1(new_n1001_), .A2(KEYINPUT119), .ZN(new_n1002_));
  NAND2_X1  g801(.A1(new_n1001_), .A2(KEYINPUT119), .ZN(new_n1003_));
  XNOR2_X1  g802(.A(KEYINPUT61), .B(G155gat), .ZN(new_n1004_));
  AND3_X1   g803(.A1(new_n1002_), .A2(new_n1003_), .A3(new_n1004_), .ZN(new_n1005_));
  AOI21_X1  g804(.A(new_n1004_), .B1(new_n1002_), .B2(new_n1003_), .ZN(new_n1006_));
  NOR2_X1   g805(.A1(new_n1005_), .A2(new_n1006_), .ZN(G1346gat));
  NAND4_X1  g806(.A1(new_n968_), .A2(new_n726_), .A3(new_n411_), .A4(new_n994_), .ZN(new_n1008_));
  NAND2_X1  g807(.A1(new_n1008_), .A2(G162gat), .ZN(new_n1009_));
  NAND2_X1  g808(.A1(new_n739_), .A2(new_n544_), .ZN(new_n1010_));
  OAI21_X1  g809(.A(new_n1009_), .B1(new_n997_), .B2(new_n1010_), .ZN(new_n1011_));
  INV_X1    g810(.A(KEYINPUT120), .ZN(new_n1012_));
  XNOR2_X1  g811(.A(new_n1011_), .B(new_n1012_), .ZN(G1347gat));
  NOR4_X1   g812(.A1(new_n821_), .A2(new_n577_), .A3(new_n607_), .A4(new_n411_), .ZN(new_n1014_));
  NAND3_X1  g813(.A1(new_n968_), .A2(new_n737_), .A3(new_n1014_), .ZN(new_n1015_));
  NAND2_X1  g814(.A1(new_n1015_), .A2(G169gat), .ZN(new_n1016_));
  NAND2_X1  g815(.A1(new_n1016_), .A2(KEYINPUT121), .ZN(new_n1017_));
  INV_X1    g816(.A(KEYINPUT121), .ZN(new_n1018_));
  NAND3_X1  g817(.A1(new_n1015_), .A2(new_n1018_), .A3(G169gat), .ZN(new_n1019_));
  NAND2_X1  g818(.A1(new_n1017_), .A2(new_n1019_), .ZN(new_n1020_));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1021_));
  NAND2_X1  g820(.A1(new_n1020_), .A2(new_n1021_), .ZN(new_n1022_));
  NAND3_X1  g821(.A1(new_n1017_), .A2(KEYINPUT62), .A3(new_n1019_), .ZN(new_n1023_));
  NAND2_X1  g822(.A1(new_n968_), .A2(new_n1014_), .ZN(new_n1024_));
  INV_X1    g823(.A(new_n1024_), .ZN(new_n1025_));
  NAND3_X1  g824(.A1(new_n1025_), .A2(new_n737_), .A3(new_n369_), .ZN(new_n1026_));
  NAND3_X1  g825(.A1(new_n1022_), .A2(new_n1023_), .A3(new_n1026_), .ZN(G1348gat));
  NAND2_X1  g826(.A1(new_n1025_), .A2(new_n291_), .ZN(new_n1028_));
  NOR2_X1   g827(.A1(new_n1028_), .A2(new_n355_), .ZN(new_n1029_));
  AOI21_X1  g828(.A(new_n1029_), .B1(new_n368_), .B2(new_n1028_), .ZN(G1349gat));
  NOR2_X1   g829(.A1(new_n1024_), .A2(new_n696_), .ZN(new_n1031_));
  MUX2_X1   g830(.A(G183gat), .B(new_n340_), .S(new_n1031_), .Z(G1350gat));
  OAI21_X1  g831(.A(G190gat), .B1(new_n1024_), .B2(new_n725_), .ZN(new_n1033_));
  NAND2_X1  g832(.A1(new_n739_), .A2(new_n343_), .ZN(new_n1034_));
  XOR2_X1   g833(.A(new_n1034_), .B(KEYINPUT122), .Z(new_n1035_));
  INV_X1    g834(.A(new_n1035_), .ZN(new_n1036_));
  OAI21_X1  g835(.A(new_n1033_), .B1(new_n1024_), .B2(new_n1036_), .ZN(new_n1037_));
  XNOR2_X1  g836(.A(new_n1037_), .B(KEYINPUT123), .ZN(G1351gat));
  NOR2_X1   g837(.A1(new_n821_), .A2(new_n653_), .ZN(new_n1039_));
  NAND2_X1  g838(.A1(new_n993_), .A2(new_n1039_), .ZN(new_n1040_));
  NOR2_X1   g839(.A1(new_n1040_), .A2(new_n339_), .ZN(new_n1041_));
  XNOR2_X1  g840(.A(KEYINPUT124), .B(G197gat), .ZN(new_n1042_));
  NOR2_X1   g841(.A1(new_n1041_), .A2(new_n1042_), .ZN(new_n1043_));
  NAND2_X1  g842(.A1(new_n447_), .A2(KEYINPUT124), .ZN(new_n1044_));
  AOI21_X1  g843(.A(new_n1043_), .B1(new_n1041_), .B2(new_n1044_), .ZN(G1352gat));
  OAI21_X1  g844(.A(KEYINPUT126), .B1(new_n449_), .B2(KEYINPUT125), .ZN(new_n1046_));
  OAI21_X1  g845(.A(new_n1046_), .B1(KEYINPUT126), .B2(new_n449_), .ZN(new_n1047_));
  NAND3_X1  g846(.A1(new_n993_), .A2(new_n291_), .A3(new_n1039_), .ZN(new_n1048_));
  MUX2_X1   g847(.A(new_n1047_), .B(new_n1046_), .S(new_n1048_), .Z(G1353gat));
  NAND3_X1  g848(.A1(new_n993_), .A2(new_n695_), .A3(new_n1039_), .ZN(new_n1050_));
  NOR2_X1   g849(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1051_));
  AND2_X1   g850(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1052_));
  NOR3_X1   g851(.A1(new_n1050_), .A2(new_n1051_), .A3(new_n1052_), .ZN(new_n1053_));
  AOI21_X1  g852(.A(new_n1053_), .B1(new_n1050_), .B2(new_n1051_), .ZN(G1354gat));
  OAI21_X1  g853(.A(G218gat), .B1(new_n1040_), .B2(new_n725_), .ZN(new_n1055_));
  NAND2_X1  g854(.A1(new_n739_), .A2(new_n454_), .ZN(new_n1056_));
  OAI21_X1  g855(.A(new_n1055_), .B1(new_n1040_), .B2(new_n1056_), .ZN(G1355gat));
endmodule


