//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT85), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G169gat), .B(G197gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT81), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n208_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n208_), .B1(new_n207_), .B2(new_n211_), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n213_), .A2(KEYINPUT82), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT82), .B1(new_n213_), .B2(new_n214_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G1gat), .B(G8gat), .Z(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n215_), .A2(new_n218_), .A3(new_n216_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G29gat), .B(G36gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT75), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n224_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G43gat), .B(G50gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n227_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n230_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT15), .A3(new_n228_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n231_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n220_), .A2(new_n221_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n239_), .B1(new_n232_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n206_), .B1(new_n241_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n239_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n243_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n242_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n240_), .A3(new_n205_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n252_), .A2(KEYINPUT86), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(KEYINPUT86), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT90), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT23), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT23), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n259_), .B(new_n261_), .C1(G183gat), .C2(G190gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT92), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT22), .B(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT91), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT89), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(KEYINPUT91), .B2(new_n268_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n264_), .A2(new_n265_), .A3(new_n269_), .A4(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G190gat), .ZN(new_n274_));
  INV_X1    g073(.A(G183gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT25), .B1(new_n275_), .B2(KEYINPUT87), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(KEYINPUT25), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n274_), .B(new_n276_), .C1(new_n277_), .C2(KEYINPUT87), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n278_), .B(KEYINPUT88), .Z(new_n279_));
  MUX2_X1   g078(.A(new_n256_), .B(new_n258_), .S(new_n260_), .Z(new_n280_));
  NOR3_X1   g079(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n271_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n281_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n279_), .A2(new_n280_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n273_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G71gat), .B(G99gat), .ZN(new_n288_));
  INV_X1    g087(.A(G43gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT30), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G227gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(G15gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n291_), .B(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n287_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT93), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n287_), .A2(new_n295_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT31), .ZN(new_n300_));
  XOR2_X1   g099(.A(G127gat), .B(G134gat), .Z(new_n301_));
  XOR2_X1   g100(.A(G113gat), .B(G120gat), .Z(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n296_), .A2(new_n297_), .A3(new_n304_), .A4(new_n298_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n300_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n303_), .B1(new_n300_), .B2(new_n305_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G155gat), .B(G162gat), .Z(new_n310_));
  OR3_X1    g109(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT94), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n311_), .B(new_n312_), .C1(new_n315_), .C2(KEYINPUT2), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n315_), .A2(KEYINPUT2), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n310_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n310_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G141gat), .ZN(new_n321_));
  INV_X1    g120(.A(G148gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n320_), .A2(new_n313_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n326_), .A2(new_n303_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n303_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n327_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n331_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G85gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT0), .B(G57gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n331_), .B(new_n343_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT27), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT25), .B(G183gat), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n274_), .A2(new_n348_), .B1(new_n284_), .B2(new_n270_), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT98), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n259_), .A2(new_n261_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(new_n281_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G211gat), .B(G218gat), .Z(new_n354_));
  INV_X1    g153(.A(G197gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G204gat), .ZN(new_n356_));
  INV_X1    g155(.A(G204gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G197gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(KEYINPUT21), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT96), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n359_), .A2(KEYINPUT21), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n362_), .A2(new_n354_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n356_), .A2(new_n358_), .A3(KEYINPUT95), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n364_), .B(KEYINPUT21), .C1(KEYINPUT95), .C2(new_n356_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n280_), .B1(G183gat), .B2(G190gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n282_), .A3(new_n268_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n353_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT99), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n361_), .A2(new_n366_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n287_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n371_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n378_), .A2(KEYINPUT20), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .A4(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n273_), .A2(new_n367_), .A3(new_n286_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n353_), .A2(new_n369_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n373_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n383_), .A3(KEYINPUT20), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n377_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT18), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  AND3_X1   g188(.A1(new_n380_), .A2(new_n385_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n347_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n326_), .A2(KEYINPUT29), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n373_), .A2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n395_), .A2(G228gat), .A3(G233gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(G228gat), .B2(G233gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n393_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT97), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n326_), .A2(KEYINPUT29), .ZN(new_n400_));
  XOR2_X1   g199(.A(G22gat), .B(G50gat), .Z(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT28), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n400_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  OR3_X1    g203(.A1(new_n396_), .A2(new_n397_), .A3(new_n393_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n398_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n399_), .A2(new_n405_), .A3(new_n398_), .A4(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n380_), .A2(new_n385_), .A3(new_n389_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n384_), .A2(new_n377_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n370_), .A2(KEYINPUT20), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n378_), .B1(new_n412_), .B2(new_n374_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(KEYINPUT27), .B(new_n410_), .C1(new_n414_), .C2(new_n389_), .ZN(new_n415_));
  AND4_X1   g214(.A1(new_n346_), .A2(new_n392_), .A3(new_n409_), .A4(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n391_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n344_), .A2(KEYINPUT100), .ZN(new_n418_));
  INV_X1    g217(.A(new_n336_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n330_), .A3(new_n333_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n343_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n418_), .A2(KEYINPUT33), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n418_), .A2(KEYINPUT33), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n417_), .A2(new_n422_), .A3(new_n410_), .A4(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n389_), .A2(KEYINPUT32), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n380_), .A2(new_n385_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n426_), .B(new_n345_), .C1(new_n425_), .C2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n409_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n309_), .B1(new_n416_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n409_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n306_), .A2(new_n307_), .A3(new_n345_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT101), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n392_), .A2(new_n433_), .A3(new_n415_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n392_), .B2(new_n415_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n431_), .B(new_n432_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n255_), .B1(new_n430_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G120gat), .B(G148gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT5), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G176gat), .B(G204gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G64gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G71gat), .B(G78gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT11), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(KEYINPUT11), .ZN(new_n446_));
  INV_X1    g245(.A(new_n444_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n443_), .A2(KEYINPUT11), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n445_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G99gat), .A2(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT6), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(G99gat), .A3(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  OR3_X1    g255(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT65), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n456_), .A2(new_n457_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n464_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G85gat), .ZN(new_n469_));
  INV_X1    g268(.A(G92gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT66), .A3(new_n465_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n462_), .A2(new_n463_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n463_), .B1(new_n462_), .B2(new_n473_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT64), .B(G92gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT9), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(G85gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(KEYINPUT9), .A3(new_n465_), .ZN(new_n480_));
  OR2_X1    g279(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n481_));
  INV_X1    g280(.A(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n479_), .A2(new_n456_), .A3(new_n480_), .A4(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n451_), .B1(new_n476_), .B2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(KEYINPUT12), .B(new_n445_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n485_), .A2(KEYINPUT68), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n456_), .A2(new_n480_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n484_), .A4(new_n479_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n492_), .B1(new_n476_), .B2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n485_), .B(new_n450_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT70), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G230gat), .A2(G233gat), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n490_), .B(new_n498_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(KEYINPUT67), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n462_), .A2(new_n473_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT8), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n462_), .A2(new_n463_), .A3(new_n473_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT67), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n485_), .A4(new_n450_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n505_), .A2(new_n487_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n501_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n442_), .B1(new_n504_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n504_), .A2(new_n514_), .A3(new_n442_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT72), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT13), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(KEYINPUT13), .A3(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT73), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT79), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n476_), .A2(new_n486_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT35), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G232gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n532_), .A2(new_n231_), .B1(new_n533_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT77), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n537_), .A2(new_n533_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n509_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT76), .B1(new_n237_), .B2(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n237_), .A2(new_n543_), .A3(KEYINPUT76), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n542_), .B(new_n538_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n538_), .B1(new_n545_), .B2(new_n544_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT78), .ZN(new_n551_));
  XOR2_X1   g350(.A(G134gat), .B(G162gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n531_), .B1(new_n549_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n546_), .A2(new_n548_), .A3(KEYINPUT79), .A4(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n553_), .B(KEYINPUT36), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n549_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n561_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n549_), .B2(KEYINPUT80), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT80), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n546_), .A2(new_n548_), .A3(new_n566_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n556_), .A2(new_n558_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n563_), .B1(new_n568_), .B2(KEYINPUT37), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n222_), .A2(new_n451_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n220_), .A2(new_n221_), .A3(new_n450_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT83), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n572_), .B(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G127gat), .B(G155gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n576_), .A2(KEYINPUT17), .A3(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n581_), .B(KEYINPUT17), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n582_), .B1(new_n576_), .B2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n569_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n437_), .A2(new_n530_), .A3(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n345_), .B(KEYINPUT102), .Z(new_n588_));
  NOR3_X1   g387(.A1(new_n587_), .A2(G1gat), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT38), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT103), .Z(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n568_), .B1(new_n430_), .B2(new_n436_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n526_), .A2(new_n251_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(new_n585_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT104), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n345_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n592_), .B1(new_n598_), .B2(G1gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n591_), .B1(new_n599_), .B2(new_n589_), .ZN(G1324gat));
  INV_X1    g399(.A(new_n587_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n434_), .A2(new_n435_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(new_n210_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  INV_X1    g404(.A(new_n596_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n603_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n605_), .B1(new_n607_), .B2(G8gat), .ZN(new_n608_));
  AOI211_X1 g407(.A(KEYINPUT39), .B(new_n210_), .C1(new_n606_), .C2(new_n603_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n604_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g410(.A1(new_n601_), .A2(new_n293_), .A3(new_n308_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n597_), .A2(new_n308_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n613_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT41), .B1(new_n613_), .B2(G15gat), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(G1326gat));
  OR3_X1    g415(.A1(new_n587_), .A2(G22gat), .A3(new_n431_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n597_), .A2(new_n409_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n619_));
  AND3_X1   g418(.A1(new_n618_), .A2(G22gat), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n618_), .B2(G22gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n620_), .B2(new_n621_), .ZN(G1327gat));
  NAND2_X1  g421(.A1(new_n565_), .A2(new_n567_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n559_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n585_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n525_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n437_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n345_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n430_), .A2(new_n436_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n569_), .A3(new_n631_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n624_), .A2(new_n560_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n430_), .B2(new_n436_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n631_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n632_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n594_), .A2(new_n625_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(KEYINPUT44), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT44), .B1(new_n638_), .B2(new_n639_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n588_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(G29gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n629_), .B1(new_n643_), .B2(new_n645_), .ZN(G1328gat));
  INV_X1    g445(.A(G36gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n628_), .A2(new_n647_), .A3(new_n603_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT45), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n641_), .A2(new_n602_), .A3(new_n642_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(new_n647_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT46), .B(new_n649_), .C1(new_n650_), .C2(new_n647_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  NOR2_X1   g454(.A1(new_n309_), .A2(new_n289_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n643_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n289_), .B1(new_n627_), .B2(new_n309_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT47), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT47), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n657_), .A2(new_n661_), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1330gat));
  AOI21_X1  g462(.A(G50gat), .B1(new_n628_), .B2(new_n409_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n409_), .A2(G50gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n643_), .B2(new_n665_), .ZN(G1331gat));
  NAND2_X1  g465(.A1(new_n630_), .A2(new_n252_), .ZN(new_n667_));
  NOR4_X1   g466(.A1(new_n667_), .A2(new_n585_), .A3(new_n526_), .A4(new_n569_), .ZN(new_n668_));
  INV_X1    g467(.A(G57gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n644_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n530_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n585_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n593_), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G57gat), .B1(new_n673_), .B2(new_n346_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n674_), .ZN(G1332gat));
  INV_X1    g474(.A(G64gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n668_), .A2(new_n676_), .A3(new_n603_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n673_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n676_), .B1(new_n678_), .B2(new_n603_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n680_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n683_));
  AND3_X1   g482(.A1(new_n681_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n677_), .B1(new_n684_), .B2(new_n685_), .ZN(G1333gat));
  INV_X1    g485(.A(G71gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n668_), .A2(new_n687_), .A3(new_n308_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n678_), .B2(new_n308_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n689_), .A2(new_n690_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(G1334gat));
  OAI21_X1  g492(.A(G78gat), .B1(new_n673_), .B2(new_n431_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT50), .ZN(new_n695_));
  INV_X1    g494(.A(G78gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n668_), .A2(new_n696_), .A3(new_n409_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1335gat));
  NAND3_X1  g497(.A1(new_n671_), .A2(new_n568_), .A3(new_n585_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT110), .B1(new_n699_), .B2(new_n667_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n530_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n667_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n702_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n469_), .B(new_n644_), .C1(new_n701_), .C2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n525_), .A2(new_n585_), .A3(new_n252_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n638_), .A2(KEYINPUT111), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n632_), .B(new_n710_), .C1(new_n634_), .C2(new_n637_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n345_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n707_), .B1(new_n713_), .B2(new_n469_), .ZN(G1336gat));
  OAI21_X1  g513(.A(new_n603_), .B1(new_n701_), .B2(new_n706_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n603_), .A2(new_n477_), .ZN(new_n716_));
  AOI22_X1  g515(.A1(new_n715_), .A2(new_n470_), .B1(new_n712_), .B2(new_n716_), .ZN(G1337gat));
  AND2_X1   g516(.A1(new_n481_), .A2(new_n483_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n308_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n700_), .B2(new_n705_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n709_), .A2(new_n711_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n708_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n308_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n720_), .B1(new_n723_), .B2(G99gat), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n725_), .ZN(new_n727_));
  AOI211_X1 g526(.A(new_n727_), .B(new_n720_), .C1(new_n723_), .C2(G99gat), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1338gat));
  OAI211_X1 g528(.A(new_n482_), .B(new_n409_), .C1(new_n701_), .C2(new_n706_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n482_), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n708_), .A2(new_n431_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n638_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n730_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT53), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n730_), .B(new_n741_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1339gat));
  NAND2_X1  g542(.A1(new_n526_), .A2(new_n672_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT54), .B1(new_n744_), .B2(new_n569_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT54), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n633_), .A2(new_n746_), .A3(new_n526_), .A4(new_n672_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n520_), .A2(new_n251_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n502_), .A2(new_n503_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n450_), .B1(new_n509_), .B2(new_n485_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n498_), .B1(new_n753_), .B2(new_n488_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OR3_X1    g556(.A1(new_n752_), .A2(new_n751_), .A3(new_n754_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759_));
  INV_X1    g558(.A(new_n499_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n754_), .B2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n490_), .A2(KEYINPUT115), .A3(new_n499_), .A4(new_n498_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n513_), .A3(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n504_), .A2(KEYINPUT114), .A3(new_n751_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n757_), .A2(new_n758_), .A3(new_n763_), .A4(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n441_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n441_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n750_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT116), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n750_), .B(new_n770_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n239_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n232_), .A2(new_n238_), .A3(new_n246_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n206_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n250_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n771_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n624_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n568_), .A2(new_n781_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n520_), .A2(new_n251_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n765_), .A2(new_n441_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n441_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n778_), .B1(new_n789_), .B2(new_n770_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n771_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n783_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n520_), .A2(new_n795_), .A3(new_n775_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n520_), .B2(new_n775_), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n796_), .A2(new_n797_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI221_X1 g599(.A(KEYINPUT58), .B1(new_n766_), .B2(new_n767_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n569_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n779_), .A2(KEYINPUT118), .A3(new_n783_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n782_), .A2(new_n794_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n749_), .B1(new_n804_), .B2(new_n585_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n602_), .A2(new_n431_), .A3(new_n308_), .A4(new_n644_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G113gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n251_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n255_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n813_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n526_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n807_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n530_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n815_), .ZN(G1341gat));
  AOI21_X1  g618(.A(G127gat), .B1(new_n807_), .B2(new_n625_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n810_), .A2(new_n812_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(G127gat), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n625_), .A2(KEYINPUT119), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(G127gat), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n820_), .B1(new_n821_), .B2(new_n825_), .ZN(G1342gat));
  AOI21_X1  g625(.A(new_n777_), .B1(new_n768_), .B2(KEYINPUT116), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n568_), .B1(new_n827_), .B2(new_n771_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n802_), .B1(new_n828_), .B2(KEYINPUT57), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n779_), .A2(KEYINPUT118), .A3(new_n783_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT118), .B1(new_n779_), .B2(new_n783_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n748_), .B1(new_n832_), .B2(new_n625_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n806_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n568_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(G134gat), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n835_), .A2(KEYINPUT120), .A3(new_n836_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n633_), .A2(new_n836_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n839_), .A2(new_n840_), .B1(new_n821_), .B2(new_n841_), .ZN(G1343gat));
  XNOR2_X1  g641(.A(KEYINPUT121), .B(G141gat), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n602_), .A2(new_n409_), .A3(new_n309_), .A4(new_n644_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n805_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n847_), .B2(new_n251_), .ZN(new_n848_));
  NOR4_X1   g647(.A1(new_n805_), .A2(KEYINPUT122), .A3(new_n252_), .A4(new_n846_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n844_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n846_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n833_), .A2(new_n251_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT122), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n847_), .A2(new_n845_), .A3(new_n251_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n843_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n850_), .A2(new_n855_), .ZN(G1344gat));
  NAND2_X1  g655(.A1(new_n847_), .A2(new_n671_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g657(.A1(new_n830_), .A2(new_n831_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n829_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n625_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n625_), .B(new_n851_), .C1(new_n861_), .C2(new_n749_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT123), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n833_), .A2(new_n864_), .A3(new_n625_), .A4(new_n851_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n863_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1346gat));
  INV_X1    g668(.A(G162gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n847_), .A2(new_n870_), .A3(new_n568_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n805_), .A2(new_n633_), .A3(new_n846_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n870_), .B2(new_n872_), .ZN(G1347gat));
  NOR4_X1   g672(.A1(new_n602_), .A2(new_n409_), .A3(new_n309_), .A4(new_n644_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n833_), .A2(new_n251_), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(G169gat), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(KEYINPUT62), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(KEYINPUT124), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n874_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n805_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n266_), .A3(new_n251_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n875_), .B(new_n878_), .C1(new_n877_), .C2(KEYINPUT62), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(new_n884_), .A3(new_n885_), .ZN(G1348gat));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n267_), .A3(new_n525_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n805_), .A2(new_n530_), .A3(new_n882_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n267_), .B2(new_n888_), .ZN(G1349gat));
  NAND2_X1  g688(.A1(new_n883_), .A2(new_n625_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n348_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n275_), .B2(new_n890_), .ZN(G1350gat));
  NAND2_X1  g691(.A1(new_n883_), .A2(new_n569_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G190gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n883_), .A2(new_n274_), .A3(new_n568_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1351gat));
  NOR3_X1   g695(.A1(new_n308_), .A2(new_n431_), .A3(new_n345_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT125), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n602_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT126), .B1(new_n805_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n902_), .B(new_n899_), .C1(new_n861_), .C2(new_n749_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G197gat), .B1(new_n904_), .B2(new_n251_), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n355_), .B(new_n252_), .C1(new_n901_), .C2(new_n903_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1352gat));
  AOI21_X1  g706(.A(new_n902_), .B1(new_n833_), .B2(new_n899_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n805_), .A2(KEYINPUT126), .A3(new_n900_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n671_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G204gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n904_), .A2(new_n357_), .A3(new_n671_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1353gat));
  OR2_X1    g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n904_), .B2(new_n625_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT63), .B(G211gat), .ZN(new_n916_));
  AOI211_X1 g715(.A(new_n585_), .B(new_n916_), .C1(new_n901_), .C2(new_n903_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1354gat));
  NAND2_X1  g717(.A1(new_n904_), .A2(new_n568_), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT127), .B(G218gat), .Z(new_n920_));
  NOR2_X1   g719(.A1(new_n633_), .A2(new_n920_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n919_), .A2(new_n920_), .B1(new_n904_), .B2(new_n921_), .ZN(G1355gat));
endmodule


