//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT10), .B(G99gat), .Z(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G92gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(G85gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G85gat), .B(G92gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n207_), .B(new_n210_), .C1(new_n209_), .C2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n211_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n213_), .B1(new_n216_), .B2(new_n204_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(KEYINPUT8), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n214_), .B(KEYINPUT7), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n211_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n212_), .B1(new_n218_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G50gat), .ZN(new_n225_));
  OR2_X1    g024(.A1(G29gat), .A2(G36gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G29gat), .A2(G36gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT70), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT70), .B1(new_n226_), .B2(new_n227_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n229_), .A2(G43gat), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G43gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G29gat), .B(G36gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n232_), .B1(new_n235_), .B2(new_n228_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n225_), .B1(new_n231_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(G43gat), .B1(new_n229_), .B2(new_n230_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n232_), .A3(new_n228_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(G50gat), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n224_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT15), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n237_), .A2(KEYINPUT15), .A3(new_n240_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n242_), .B1(new_n246_), .B2(new_n224_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G232gat), .A2(G233gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT34), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT35), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n252_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n251_), .A2(KEYINPUT35), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n249_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G190gat), .B(G218gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G134gat), .ZN(new_n258_));
  INV_X1    g057(.A(G162gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT36), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n245_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT15), .B1(new_n237_), .B2(new_n240_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n224_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n242_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n253_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n251_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n265_), .A2(new_n248_), .A3(new_n266_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n255_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n256_), .A2(new_n262_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n260_), .A2(new_n261_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n256_), .B2(new_n271_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G127gat), .B(G134gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G113gat), .B(G120gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT87), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT86), .B(G15gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G71gat), .B(G99gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n291_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G227gat), .A2(G233gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT85), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT31), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(new_n232_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  INV_X1    g098(.A(G176gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT81), .B1(new_n301_), .B2(G169gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT22), .B(G169gat), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n300_), .B(new_n302_), .C1(new_n303_), .C2(KEYINPUT81), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT23), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(G183gat), .A3(G190gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT82), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n307_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(G183gat), .ZN(new_n312_));
  AND2_X1   g111(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n316_), .A2(KEYINPUT83), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(KEYINPUT83), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n299_), .B(new_n304_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n306_), .A2(new_n308_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n321_));
  INV_X1    g120(.A(G169gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n300_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT24), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT78), .B(G190gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT26), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(KEYINPUT25), .B(G183gat), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n331_), .A2(KEYINPUT79), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT79), .B1(new_n331_), .B2(new_n333_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n320_), .B(new_n327_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n323_), .A2(KEYINPUT24), .A3(new_n299_), .A4(new_n324_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n319_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n298_), .A2(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n298_), .A2(new_n339_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n294_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n340_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n293_), .A3(new_n292_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n347_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(G155gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n259_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G141gat), .B(G148gat), .Z(new_n358_));
  NAND2_X1  g157(.A1(new_n346_), .A2(KEYINPUT1), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT88), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n346_), .A2(KEYINPUT1), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT88), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n346_), .A2(new_n362_), .A3(KEYINPUT1), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .A4(new_n357_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n355_), .A2(new_n357_), .B1(new_n358_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT28), .Z(new_n368_));
  AND2_X1   g167(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(G204gat), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT21), .ZN(new_n372_));
  INV_X1    g171(.A(G197gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(G204gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT90), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n373_), .ZN(new_n380_));
  INV_X1    g179(.A(G204gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT91), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n373_), .A2(G204gat), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n380_), .A2(KEYINPUT91), .A3(new_n381_), .A4(new_n382_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n378_), .B1(KEYINPUT21), .B2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n371_), .A2(new_n375_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n390_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT94), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(KEYINPUT21), .ZN(new_n393_));
  INV_X1    g192(.A(new_n378_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT94), .ZN(new_n396_));
  INV_X1    g195(.A(new_n391_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n350_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n354_), .A2(new_n348_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n346_), .A3(new_n357_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n364_), .A2(new_n358_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n392_), .A2(new_n398_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G228gat), .ZN(new_n407_));
  INV_X1    g206(.A(G233gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n403_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n409_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT92), .B1(new_n395_), .B2(new_n397_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n389_), .A2(new_n417_), .A3(new_n391_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n414_), .B(new_n415_), .C1(new_n416_), .C2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G22gat), .B(G50gat), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n410_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n410_), .B2(new_n419_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n368_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n410_), .A2(new_n419_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n420_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n368_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n410_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n423_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n423_), .B2(new_n429_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n345_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n430_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n421_), .A2(new_n422_), .A3(new_n368_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n427_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n345_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n423_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n433_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT103), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G8gat), .B(G36gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G64gat), .B(G92gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT95), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n310_), .A2(new_n311_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT24), .B1(new_n323_), .B2(new_n324_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n327_), .A2(KEYINPUT95), .A3(new_n311_), .A4(new_n310_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT26), .B(G190gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n333_), .A2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n452_), .A2(new_n453_), .A3(new_n337_), .A4(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n320_), .B1(G183gat), .B2(G190gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n299_), .B(KEYINPUT96), .Z(new_n458_));
  INV_X1    g257(.A(new_n303_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n457_), .B(new_n458_), .C1(G176gat), .C2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n395_), .A2(new_n397_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G226gat), .A2(G233gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT19), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n463_), .A2(KEYINPUT20), .A3(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n417_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n395_), .A2(KEYINPUT92), .A3(new_n397_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n339_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT97), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n339_), .A3(KEYINPUT97), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n467_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n461_), .A2(new_n462_), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT20), .B(new_n476_), .C1(new_n470_), .C2(new_n339_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n477_), .A2(new_n465_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n448_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n463_), .A2(KEYINPUT20), .A3(new_n466_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n474_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT97), .B1(new_n470_), .B2(new_n339_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n465_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n447_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n479_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n442_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  AOI211_X1 g288(.A(KEYINPUT103), .B(new_n487_), .C1(new_n479_), .C2(new_n485_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G85gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT0), .ZN(new_n494_));
  INV_X1    g293(.A(G57gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n403_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT4), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n365_), .A2(new_n280_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT99), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT99), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n365_), .A2(new_n502_), .A3(new_n280_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n497_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n499_), .B1(new_n504_), .B2(KEYINPUT4), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G225gat), .A2(G233gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n504_), .A2(new_n506_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n496_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n507_), .B2(new_n505_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n496_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n477_), .A2(new_n465_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n392_), .A2(new_n398_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT100), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n461_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n456_), .A2(KEYINPUT100), .A3(new_n460_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT20), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT101), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT101), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n524_), .A3(KEYINPUT20), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n473_), .A2(new_n474_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n516_), .B1(new_n527_), .B2(new_n465_), .ZN(new_n528_));
  OAI211_X1 g327(.A(KEYINPUT27), .B(new_n485_), .C1(new_n528_), .C2(new_n447_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n441_), .A2(new_n491_), .A3(new_n515_), .A4(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n504_), .A2(new_n506_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT33), .B1(new_n532_), .B2(new_n496_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n510_), .ZN(new_n534_));
  OAI211_X1 g333(.A(KEYINPUT33), .B(new_n496_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n534_), .A2(new_n485_), .A3(new_n479_), .A4(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n447_), .A2(KEYINPUT32), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n528_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n483_), .A2(new_n484_), .A3(new_n537_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n514_), .A2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n536_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n431_), .A2(new_n432_), .A3(new_n438_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n277_), .B1(new_n530_), .B2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n544_), .B(KEYINPUT106), .Z(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT72), .B(G1gat), .Z(new_n546_));
  INV_X1    g345(.A(G8gat), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT14), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(G1gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(G15gat), .B(G22gat), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT72), .B(G1gat), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(G8gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(G1gat), .B1(new_n555_), .B2(new_n550_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n547_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n552_), .A2(G8gat), .A3(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT73), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n560_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G57gat), .B(G64gat), .Z(new_n564_));
  INV_X1    g363(.A(KEYINPUT11), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(G71gat), .ZN(new_n567_));
  INV_X1    g366(.A(G78gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(KEYINPUT66), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT66), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n564_), .A2(new_n565_), .B1(G71gat), .B2(G78gat), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n569_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n564_), .A2(new_n565_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n572_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(KEYINPUT66), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(new_n573_), .A3(new_n569_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n576_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n563_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G183gat), .B(G211gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT17), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n583_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n593_), .B2(new_n583_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n545_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n224_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n577_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n221_), .B(new_n222_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n579_), .A2(new_n580_), .A3(new_n576_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n212_), .A4(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT67), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT64), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n603_), .B(new_n605_), .C1(new_n602_), .C2(new_n601_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT5), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(G176gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(G204gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n597_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n605_), .ZN(new_n614_));
  OR2_X1    g413(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n224_), .B(new_n615_), .C1(new_n578_), .C2(new_n581_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n601_), .A4(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n606_), .A2(new_n610_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n610_), .B(KEYINPUT69), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n606_), .A2(new_n617_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT13), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n558_), .A2(new_n559_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n246_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G229gat), .A2(G233gat), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT76), .ZN(new_n630_));
  INV_X1    g429(.A(new_n241_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n560_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n560_), .B2(new_n631_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n628_), .B(new_n629_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT77), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(new_n322_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(new_n373_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT76), .B1(new_n627_), .B2(new_n241_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n560_), .A2(new_n631_), .A3(new_n630_), .ZN(new_n641_));
  AOI22_X1  g440(.A1(new_n640_), .A2(new_n641_), .B1(new_n241_), .B2(new_n627_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n634_), .B(new_n639_), .C1(new_n642_), .C2(new_n629_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI22_X1  g443(.A1(new_n632_), .A2(new_n633_), .B1(new_n631_), .B2(new_n560_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n629_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n639_), .B1(new_n647_), .B2(new_n634_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n626_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n596_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n515_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT37), .B1(new_n272_), .B2(new_n275_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n271_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n269_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n273_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT37), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n256_), .A2(new_n271_), .A3(new_n262_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n655_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n595_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT75), .Z(new_n664_));
  AOI21_X1  g463(.A(new_n651_), .B1(new_n530_), .B2(new_n543_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT104), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n514_), .A3(new_n546_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT105), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT38), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT38), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n654_), .B1(new_n670_), .B2(new_n671_), .ZN(G1324gat));
  NAND2_X1  g471(.A1(new_n486_), .A2(new_n488_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT103), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n486_), .A2(new_n442_), .A3(new_n488_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n529_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G8gat), .B1(new_n653_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT39), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(G8gat), .C1(new_n653_), .C2(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n667_), .A2(new_n547_), .A3(new_n676_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n682_), .A2(KEYINPUT40), .A3(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1325gat));
  OAI21_X1  g487(.A(G15gat), .B1(new_n653_), .B2(new_n345_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT41), .Z(new_n690_));
  NOR3_X1   g489(.A1(new_n666_), .A2(G15gat), .A3(new_n345_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT107), .Z(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n431_), .A2(new_n432_), .ZN(new_n694_));
  OR3_X1    g493(.A1(new_n666_), .A2(G22gat), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G22gat), .B1(new_n653_), .B2(new_n694_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT108), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n698_), .B(G22gat), .C1(new_n653_), .C2(new_n694_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n697_), .A2(KEYINPUT42), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT42), .B1(new_n697_), .B2(new_n699_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n695_), .B1(new_n700_), .B2(new_n701_), .ZN(G1327gat));
  NOR2_X1   g501(.A1(new_n651_), .A2(new_n594_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n272_), .A2(new_n275_), .A3(KEYINPUT37), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n659_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI211_X1 g505(.A(KEYINPUT43), .B(new_n706_), .C1(new_n530_), .C2(new_n543_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n431_), .A2(new_n432_), .A3(new_n345_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n438_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n515_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n543_), .B1(new_n711_), .B2(new_n676_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n708_), .B1(new_n712_), .B2(new_n662_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n703_), .B1(new_n707_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT44), .B(new_n703_), .C1(new_n707_), .C2(new_n713_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n514_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT109), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n716_), .A2(new_n720_), .A3(new_n514_), .A4(new_n717_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(G29gat), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n719_), .A2(KEYINPUT110), .A3(G29gat), .A4(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n276_), .A2(new_n594_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n665_), .A2(new_n727_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n728_), .A2(G29gat), .A3(new_n515_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT111), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n726_), .A2(new_n732_), .A3(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1328gat));
  NOR3_X1   g533(.A1(new_n728_), .A2(G36gat), .A3(new_n677_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT45), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n716_), .A2(new_n676_), .A3(new_n717_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G36gat), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT46), .ZN(G1329gat));
  NAND3_X1  g538(.A1(new_n716_), .A2(new_n438_), .A3(new_n717_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G43gat), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n728_), .A2(G43gat), .A3(new_n345_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT112), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g545(.A(new_n694_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n716_), .A2(new_n747_), .A3(new_n717_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n225_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT113), .ZN(new_n750_));
  OAI22_X1  g549(.A1(new_n748_), .A2(new_n225_), .B1(new_n728_), .B2(new_n750_), .ZN(G1331gat));
  NOR2_X1   g550(.A1(new_n626_), .A2(new_n650_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n596_), .A2(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n753_), .A2(new_n495_), .A3(new_n515_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT114), .Z(new_n755_));
  AND2_X1   g554(.A1(new_n712_), .A2(new_n752_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n664_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n514_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1332gat));
  OAI21_X1  g558(.A(G64gat), .B1(new_n753_), .B2(new_n677_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(G64gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n757_), .A2(new_n763_), .A3(new_n676_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n753_), .B2(new_n345_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT49), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(G71gat), .C1(new_n753_), .C2(new_n345_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n757_), .A2(new_n567_), .A3(new_n438_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT116), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n774_), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1334gat));
  OAI21_X1  g575(.A(G78gat), .B1(new_n753_), .B2(new_n694_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT50), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n757_), .A2(new_n568_), .A3(new_n747_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1335gat));
  AND2_X1   g579(.A1(new_n756_), .A2(new_n727_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n514_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n707_), .A2(new_n713_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n595_), .A3(new_n752_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT117), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n514_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n782_), .B1(new_n786_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g586(.A(G92gat), .B1(new_n781_), .B2(new_n676_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n785_), .A2(new_n676_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n208_), .ZN(G1337gat));
  NAND3_X1  g589(.A1(new_n781_), .A2(new_n206_), .A3(new_n438_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n783_), .A2(new_n595_), .A3(new_n438_), .A4(new_n752_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n792_), .A2(KEYINPUT118), .A3(G99gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT118), .B1(new_n792_), .B2(G99gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT119), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n791_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n796_), .A2(KEYINPUT51), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n796_), .B2(new_n798_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1338gat));
  NAND3_X1  g600(.A1(new_n781_), .A2(new_n205_), .A3(new_n747_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n784_), .A2(new_n694_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G106gat), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(KEYINPUT52), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(KEYINPUT52), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT53), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(new_n802_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1339gat));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n598_), .A2(new_n600_), .B1(new_n599_), .B2(new_n212_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n616_), .B(new_n601_), .C1(new_n813_), .C2(new_n611_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n814_), .B2(new_n605_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n605_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n814_), .A2(new_n812_), .A3(new_n605_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n620_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT56), .B(new_n620_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n628_), .B(new_n646_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n638_), .B(new_n824_), .C1(new_n642_), .C2(new_n646_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n643_), .A2(new_n825_), .A3(new_n618_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT120), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n643_), .A2(new_n825_), .A3(new_n828_), .A4(new_n618_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT58), .B1(new_n823_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT121), .B1(new_n831_), .B2(new_n706_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n821_), .A2(new_n822_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT58), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n835_), .B(new_n662_), .C1(new_n833_), .C2(KEYINPUT58), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n832_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n618_), .B1(new_n644_), .B2(new_n648_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n643_), .A2(new_n825_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n622_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n843_), .B2(new_n277_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT57), .B(new_n276_), .C1(new_n840_), .C2(new_n842_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n595_), .B1(new_n837_), .B2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n706_), .A2(new_n649_), .A3(new_n594_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n626_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT54), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n663_), .A2(new_n851_), .A3(new_n649_), .A4(new_n626_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n847_), .A2(KEYINPUT122), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  INV_X1    g654(.A(new_n839_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n814_), .A2(new_n605_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT55), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n617_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n818_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT56), .B1(new_n861_), .B2(new_n620_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n822_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n856_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n842_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n866_), .B2(new_n276_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n845_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n832_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n594_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n853_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n855_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n854_), .A2(new_n873_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n676_), .A2(new_n515_), .A3(new_n440_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877_), .B2(new_n650_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT59), .B1(new_n847_), .B2(new_n853_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n876_), .A2(KEYINPUT59), .B1(new_n875_), .B2(new_n879_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n650_), .A2(G113gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n878_), .B1(new_n880_), .B2(new_n881_), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n626_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n877_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n883_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n880_), .A2(new_n849_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n883_), .ZN(G1341gat));
  AOI21_X1  g686(.A(G127gat), .B1(new_n877_), .B2(new_n594_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n594_), .A2(G127gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n880_), .B2(new_n889_), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(new_n877_), .B2(new_n277_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n662_), .A2(G134gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT123), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n880_), .B2(new_n893_), .ZN(G1343gat));
  NOR2_X1   g693(.A1(new_n676_), .A2(new_n515_), .ZN(new_n895_));
  AND4_X1   g694(.A1(new_n710_), .A2(new_n854_), .A3(new_n873_), .A4(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n650_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n849_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G148gat), .ZN(G1345gat));
  AND3_X1   g699(.A1(new_n854_), .A2(new_n873_), .A3(new_n710_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n594_), .A4(new_n895_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n854_), .A2(new_n873_), .A3(new_n710_), .A4(new_n895_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT124), .B1(new_n905_), .B2(new_n595_), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n903_), .A2(new_n904_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n904_), .B1(new_n903_), .B2(new_n906_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n356_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n902_), .B1(new_n896_), .B2(new_n594_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n905_), .A2(KEYINPUT124), .A3(new_n595_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT61), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n903_), .A2(new_n904_), .A3(new_n906_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G155gat), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n909_), .A2(new_n914_), .ZN(G1346gat));
  AOI21_X1  g714(.A(G162gat), .B1(new_n896_), .B2(new_n277_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n905_), .A2(new_n259_), .A3(new_n706_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1347gat));
  AOI21_X1  g717(.A(new_n747_), .B1(new_n847_), .B2(new_n853_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n676_), .A2(new_n515_), .A3(new_n438_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT125), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n322_), .B1(new_n923_), .B2(new_n650_), .ZN(new_n924_));
  OR2_X1    g723(.A1(new_n924_), .A2(KEYINPUT62), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n650_), .A3(new_n303_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(KEYINPUT62), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(G1348gat));
  OAI21_X1  g727(.A(new_n300_), .B1(new_n922_), .B2(new_n626_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT126), .Z(new_n930_));
  AND2_X1   g729(.A1(new_n874_), .A2(new_n694_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n921_), .A2(G176gat), .A3(new_n849_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  AND2_X1   g732(.A1(new_n921_), .A2(new_n594_), .ZN(new_n934_));
  AOI21_X1  g733(.A(G183gat), .B1(new_n931_), .B2(new_n934_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n934_), .A2(new_n332_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n919_), .B2(new_n936_), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n922_), .B2(new_n706_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n277_), .A2(new_n454_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n922_), .B2(new_n939_), .ZN(G1351gat));
  AND2_X1   g739(.A1(new_n874_), .A2(new_n676_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n433_), .A2(new_n514_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT127), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n649_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n373_), .ZN(G1352gat));
  NOR2_X1   g745(.A1(new_n944_), .A2(new_n626_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(new_n381_), .ZN(G1353gat));
  INV_X1    g747(.A(new_n944_), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT63), .B(G211gat), .Z(new_n950_));
  NAND3_X1  g749(.A1(new_n949_), .A2(new_n594_), .A3(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n952_), .B1(new_n944_), .B2(new_n595_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1354gat));
  AND3_X1   g753(.A1(new_n949_), .A2(G218gat), .A3(new_n662_), .ZN(new_n955_));
  AOI21_X1  g754(.A(G218gat), .B1(new_n949_), .B2(new_n277_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n955_), .A2(new_n956_), .ZN(G1355gat));
endmodule


