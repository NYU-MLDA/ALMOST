//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(KEYINPUT65), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT10), .B(G99gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n205_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(KEYINPUT9), .A3(new_n216_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n209_), .A2(new_n210_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT8), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n219_), .A2(KEYINPUT65), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n212_), .A2(new_n217_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n202_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n234_));
  INV_X1    g033(.A(G78gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G71gat), .ZN(new_n236_));
  INV_X1    g035(.A(G71gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G78gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(G57gat), .A2(G64gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G57gat), .A2(G64gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT66), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G57gat), .ZN(new_n243_));
  INV_X1    g042(.A(G64gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G57gat), .A2(G64gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI211_X1 g047(.A(new_n234_), .B(new_n239_), .C1(new_n242_), .C2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n234_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n242_), .A2(new_n248_), .A3(new_n234_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n239_), .A3(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n231_), .A2(new_n250_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n233_), .A2(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n242_), .A2(new_n248_), .A3(new_n234_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(new_n251_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n249_), .B1(new_n258_), .B2(new_n239_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n259_), .B(new_n231_), .C1(new_n232_), .C2(new_n202_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n220_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n254_), .A2(new_n250_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT64), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n262_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  AOI211_X1 g068(.A(KEYINPUT69), .B(new_n267_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n261_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n272_), .A3(new_n255_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n273_), .B(new_n267_), .C1(new_n272_), .C2(new_n255_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G120gat), .B(G148gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(G204gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G176gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n279_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n271_), .A2(new_n274_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT13), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(KEYINPUT13), .A3(new_n282_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G226gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT19), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT92), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G211gat), .A2(G218gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n295_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT92), .B1(new_n297_), .B2(new_n292_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G197gat), .ZN(new_n300_));
  OR3_X1    g099(.A1(new_n300_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT91), .B1(new_n300_), .B2(G204gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT89), .B(G197gat), .ZN(new_n303_));
  INV_X1    g102(.A(G204gat), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n301_), .B(new_n302_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n299_), .B1(new_n305_), .B2(KEYINPUT21), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n300_), .A2(KEYINPUT89), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G197gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n309_), .A3(new_n304_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT90), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT90), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n303_), .A2(new_n312_), .A3(new_n304_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n311_), .B(new_n313_), .C1(G197gat), .C2(new_n304_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n306_), .B1(KEYINPUT21), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G169gat), .ZN(new_n316_));
  INV_X1    g115(.A(G176gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT22), .B(G169gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(new_n317_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT95), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(KEYINPUT23), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(new_n323_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n322_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT82), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT82), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT23), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n332_), .A3(new_n323_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(KEYINPUT23), .B2(new_n323_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n327_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT95), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n321_), .B1(new_n328_), .B2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n304_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n302_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n300_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT21), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n341_), .A2(new_n299_), .A3(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n325_), .A2(new_n323_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n329_), .B1(G183gat), .B2(G190gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT24), .B1(new_n316_), .B2(new_n317_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n347_), .ZN(new_n351_));
  XOR2_X1   g150(.A(KEYINPUT26), .B(G190gat), .Z(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT25), .B(G183gat), .Z(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n346_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n355_));
  NOR4_X1   g154(.A1(new_n315_), .A2(new_n337_), .A3(new_n343_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n306_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n314_), .A2(KEYINPUT21), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n343_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT81), .B(G183gat), .ZN(new_n360_));
  OAI22_X1  g159(.A1(new_n344_), .A2(new_n345_), .B1(G190gat), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n320_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n351_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n360_), .B2(KEYINPUT25), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n363_), .B(new_n334_), .C1(new_n365_), .C2(new_n352_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n359_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n291_), .B1(new_n356_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(new_n214_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT18), .B(G64gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n373_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n359_), .A2(new_n367_), .ZN(new_n377_));
  OAI22_X1  g176(.A1(new_n315_), .A2(new_n343_), .B1(new_n337_), .B2(new_n355_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT20), .A4(new_n290_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n369_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT96), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n369_), .A2(new_n379_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n376_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n369_), .A2(KEYINPUT96), .A3(new_n376_), .A4(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n392_), .A2(new_n393_), .B1(G141gat), .B2(G148gat), .ZN(new_n394_));
  INV_X1    g193(.A(G141gat), .ZN(new_n395_));
  INV_X1    g194(.A(G148gat), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n390_), .A2(KEYINPUT1), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  OR3_X1    g197(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT2), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n392_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n398_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n398_), .A2(KEYINPUT88), .A3(new_n405_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411_));
  INV_X1    g210(.A(G50gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT28), .B(G22gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n409_), .ZN(new_n415_));
  OAI21_X1  g214(.A(G50gat), .B1(new_n415_), .B2(KEYINPUT29), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n414_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT94), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G228gat), .A2(G233gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n406_), .A2(KEYINPUT29), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n357_), .A2(new_n358_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n343_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n421_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n415_), .A2(KEYINPUT29), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(new_n427_), .A3(new_n421_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G78gat), .B(G106gat), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n428_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n420_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n422_), .B(KEYINPUT93), .ZN(new_n437_));
  OAI211_X1 g236(.A(G228gat), .B(G233gat), .C1(new_n437_), .C2(new_n359_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(new_n432_), .A3(new_n430_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n414_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n412_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n415_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n417_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n436_), .A2(new_n439_), .A3(new_n444_), .A4(KEYINPUT94), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n432_), .B1(new_n438_), .B2(new_n430_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(new_n417_), .A3(new_n443_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n435_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT101), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n376_), .B(KEYINPUT100), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n290_), .B1(new_n356_), .B2(new_n368_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT20), .A4(new_n291_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(new_n388_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n449_), .B1(new_n454_), .B2(new_n385_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n376_), .B1(new_n369_), .B2(new_n379_), .ZN(new_n456_));
  NOR4_X1   g255(.A1(new_n456_), .A2(new_n453_), .A3(KEYINPUT101), .A4(new_n388_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n389_), .B(new_n448_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT102), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n451_), .A2(new_n452_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n450_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n385_), .A2(new_n463_), .A3(KEYINPUT27), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT101), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n454_), .A2(new_n449_), .A3(new_n385_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n467_), .A2(KEYINPUT102), .A3(new_n389_), .A4(new_n448_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G120gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G113gat), .B(G120gat), .Z(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n470_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G127gat), .B(G134gat), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n469_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n473_), .A2(new_n475_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n476_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(KEYINPUT87), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n415_), .ZN(new_n487_));
  INV_X1    g286(.A(G225gat), .ZN(new_n488_));
  INV_X1    g287(.A(G233gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n479_), .A2(new_n484_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n406_), .B1(new_n483_), .B2(new_n482_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n487_), .B(new_n490_), .C1(new_n491_), .C2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(new_n485_), .B2(new_n415_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(KEYINPUT4), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G1gat), .B(G29gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(new_n213_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT0), .B(G57gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT99), .B1(new_n497_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT99), .ZN(new_n504_));
  AOI211_X1 g303(.A(new_n504_), .B(new_n501_), .C1(new_n493_), .C2(new_n496_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n493_), .A2(new_n496_), .A3(new_n501_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n503_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n362_), .A2(new_n366_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT84), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G227gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT83), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G15gat), .B(G43gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G71gat), .B(G99gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT31), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n485_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n519_), .A2(KEYINPUT31), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n519_), .A2(KEYINPUT31), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n485_), .B1(new_n525_), .B2(new_n520_), .ZN(new_n526_));
  OAI22_X1  g325(.A1(new_n524_), .A2(new_n526_), .B1(KEYINPUT84), .B2(new_n511_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n522_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n511_), .A2(KEYINPUT84), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n525_), .A2(new_n485_), .A3(new_n520_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n460_), .A2(new_n468_), .A3(new_n508_), .A4(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n389_), .B(new_n508_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n448_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n527_), .A2(new_n531_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n497_), .A2(new_n502_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n504_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n497_), .A2(KEYINPUT99), .A3(new_n502_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n506_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n384_), .A2(KEYINPUT32), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT98), .Z(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n543_), .A2(new_n383_), .B1(new_n461_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n506_), .A2(KEYINPUT97), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT33), .ZN(new_n548_));
  INV_X1    g347(.A(new_n490_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n494_), .A2(KEYINPUT4), .A3(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n550_), .B(new_n487_), .C1(new_n549_), .C2(new_n494_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n502_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n552_), .A2(new_n382_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n546_), .B(new_n448_), .C1(new_n548_), .C2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n536_), .A2(new_n537_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n288_), .B1(new_n533_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT78), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT74), .B(G1gat), .Z(new_n561_));
  INV_X1    g360(.A(G8gat), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT14), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(G22gat), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n565_), .ZN(new_n567_));
  INV_X1    g366(.A(G22gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G1gat), .B(G8gat), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n563_), .A2(new_n566_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n566_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT14), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT74), .B(G1gat), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n575_), .B2(G8gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n572_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G43gat), .B(G50gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G29gat), .B(G36gat), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n580_), .A2(new_n581_), .A3(KEYINPUT15), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G43gat), .B(G50gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n579_), .B(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT15), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n571_), .B(new_n577_), .C1(new_n582_), .C2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n577_), .A2(new_n571_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n584_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n560_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n584_), .B(KEYINPUT15), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n577_), .A2(new_n571_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT78), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n589_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n584_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n588_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n594_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n559_), .B1(new_n595_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n559_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n586_), .A2(new_n560_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n596_), .B1(new_n577_), .B2(new_n571_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n603_), .B1(new_n605_), .B2(new_n560_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n599_), .B(new_n602_), .C1(new_n606_), .C2(new_n594_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT79), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n601_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(KEYINPUT79), .B(new_n559_), .C1(new_n595_), .C2(new_n600_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT80), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(KEYINPUT80), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n556_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(G211gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT16), .B(G183gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT76), .Z(new_n622_));
  INV_X1    g421(.A(new_n619_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n622_), .A2(new_n232_), .B1(KEYINPUT17), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n264_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(new_n587_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n624_), .B(new_n628_), .C1(KEYINPUT17), .C2(new_n623_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n622_), .A2(KEYINPUT68), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT77), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT77), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n629_), .A2(new_n634_), .A3(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n590_), .A2(new_n231_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT34), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT35), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n638_), .B(new_n643_), .C1(new_n596_), .C2(new_n231_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(new_n642_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n644_), .B(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT36), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G190gat), .B(G218gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G134gat), .B(G162gat), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n649_), .B(new_n650_), .Z(new_n651_));
  XOR2_X1   g450(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n652_));
  NAND4_X1  g451(.A1(new_n647_), .A2(new_n648_), .A3(new_n651_), .A4(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n644_), .A2(new_n645_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n644_), .A2(new_n645_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n651_), .A2(new_n648_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n653_), .A2(new_n658_), .ZN(new_n659_));
  OR3_X1    g458(.A1(new_n647_), .A2(new_n648_), .A3(new_n651_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n615_), .A2(new_n637_), .A3(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n508_), .B(KEYINPUT103), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n561_), .A3(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT38), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n609_), .A2(new_n610_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n288_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n533_), .A2(new_n555_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n661_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT104), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT104), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n632_), .B(new_n673_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G1gat), .B1(new_n679_), .B2(new_n508_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n671_), .A2(new_n680_), .ZN(G1324gat));
  NAND2_X1  g480(.A1(new_n467_), .A2(new_n389_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n667_), .A2(new_n562_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n684_));
  INV_X1    g483(.A(new_n682_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n679_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n686_), .B2(G8gat), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n684_), .B(G8gat), .C1(new_n679_), .C2(new_n685_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n683_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT40), .B(new_n683_), .C1(new_n687_), .C2(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n679_), .B2(new_n537_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT41), .Z(new_n696_));
  INV_X1    g495(.A(G15gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n667_), .A2(new_n697_), .A3(new_n532_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1326gat));
  OAI21_X1  g498(.A(G22gat), .B1(new_n679_), .B2(new_n448_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT42), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(G22gat), .C1(new_n679_), .C2(new_n448_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n667_), .A2(new_n568_), .A3(new_n535_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT105), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n708_), .A3(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1327gat));
  NOR2_X1   g509(.A1(new_n636_), .A2(new_n675_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n556_), .A2(new_n614_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n713_), .B2(new_n541_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n674_), .A2(new_n666_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n674_), .A2(KEYINPUT43), .A3(new_n666_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n673_), .A3(new_n637_), .A4(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n721_), .A2(G29gat), .A3(new_n669_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT43), .B1(new_n674_), .B2(new_n666_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n666_), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n716_), .B(new_n724_), .C1(new_n533_), .C2(new_n555_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n726_), .A2(KEYINPUT44), .A3(new_n673_), .A4(new_n637_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n714_), .B1(new_n722_), .B2(new_n727_), .ZN(G1328gat));
  NOR3_X1   g527(.A1(new_n712_), .A2(G36gat), .A3(new_n685_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT45), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n721_), .A2(new_n727_), .A3(new_n682_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(G36gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n731_), .B2(G36gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n730_), .B(KEYINPUT46), .C1(new_n733_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1329gat));
  AOI21_X1  g538(.A(G43gat), .B1(new_n713_), .B2(new_n532_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT107), .Z(new_n741_));
  NAND3_X1  g540(.A1(new_n727_), .A2(G43gat), .A3(new_n532_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n721_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g544(.A1(new_n713_), .A2(new_n412_), .A3(new_n535_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n721_), .A2(new_n727_), .A3(new_n535_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n747_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT108), .B1(new_n747_), .B2(G50gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n748_), .B2(new_n749_), .ZN(G1331gat));
  AND3_X1   g549(.A1(new_n674_), .A2(KEYINPUT109), .A3(new_n672_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT109), .B1(new_n674_), .B2(new_n672_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n287_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n753_), .A2(new_n636_), .A3(new_n724_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n243_), .A3(new_n669_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n636_), .A2(new_n613_), .A3(new_n612_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n288_), .B(new_n757_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G57gat), .B1(new_n758_), .B2(new_n508_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT110), .Z(G1332gat));
  NAND3_X1  g560(.A1(new_n754_), .A2(new_n244_), .A3(new_n682_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n758_), .A2(new_n685_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(G64gat), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n763_), .B(G64gat), .C1(new_n758_), .C2(new_n685_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n762_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT111), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n762_), .B(new_n770_), .C1(new_n765_), .C2(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n758_), .B2(new_n537_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT49), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n754_), .A2(new_n237_), .A3(new_n532_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1334gat));
  OAI21_X1  g575(.A(G78gat), .B1(new_n758_), .B2(new_n448_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT50), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n754_), .A2(new_n235_), .A3(new_n535_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1335gat));
  AND2_X1   g579(.A1(new_n753_), .A2(new_n711_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n669_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n723_), .A2(new_n725_), .A3(new_n636_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n783_), .A2(new_n672_), .A3(new_n288_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n508_), .A2(new_n213_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT112), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n782_), .B1(new_n784_), .B2(new_n786_), .ZN(G1336gat));
  AOI21_X1  g586(.A(G92gat), .B1(new_n781_), .B2(new_n682_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n685_), .A2(new_n214_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n784_), .B2(new_n789_), .ZN(G1337gat));
  NAND3_X1  g589(.A1(new_n781_), .A2(new_n532_), .A3(new_n221_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n783_), .A2(new_n532_), .A3(new_n672_), .A4(new_n288_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n792_), .A2(KEYINPUT113), .A3(G99gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT113), .B1(new_n792_), .B2(G99gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n781_), .A2(new_n205_), .A3(new_n535_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n783_), .A2(new_n535_), .A3(new_n672_), .A4(new_n288_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  AND3_X1   g602(.A1(new_n460_), .A2(new_n532_), .A3(new_n468_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n669_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(KEYINPUT59), .ZN(new_n806_));
  INV_X1    g605(.A(new_n282_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n271_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n261_), .A2(new_n265_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n267_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n268_), .B1(new_n259_), .B2(new_n231_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT69), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n265_), .A2(new_n262_), .A3(new_n268_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(KEYINPUT55), .A3(new_n261_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n809_), .A2(new_n811_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n279_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n807_), .B1(new_n818_), .B2(KEYINPUT56), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n598_), .A2(new_n593_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n559_), .B(new_n820_), .C1(new_n606_), .C2(new_n593_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n822_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n823_), .A2(new_n607_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n817_), .A2(new_n826_), .A3(new_n279_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n819_), .A2(new_n825_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n819_), .A2(new_n825_), .A3(KEYINPUT58), .A4(new_n827_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n830_), .A2(new_n666_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n825_), .A2(new_n283_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n815_), .A2(KEYINPUT55), .A3(new_n261_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT55), .B1(new_n815_), .B2(new_n261_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n268_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n834_), .B(KEYINPUT56), .C1(new_n838_), .C2(new_n281_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n611_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT115), .B1(new_n817_), .B2(new_n279_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n282_), .B1(new_n841_), .B2(KEYINPUT56), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n833_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(KEYINPUT57), .A3(new_n675_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT118), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n843_), .A2(new_n846_), .A3(KEYINPUT57), .A4(new_n675_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n832_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n843_), .A2(new_n675_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n636_), .B1(new_n848_), .B2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n664_), .A2(new_n287_), .A3(new_n665_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT54), .B1(new_n756_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n756_), .A2(new_n853_), .A3(KEYINPUT54), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT114), .B(KEYINPUT54), .C1(new_n756_), .C2(new_n853_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n806_), .B1(new_n852_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n632_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n832_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n672_), .B1(new_n841_), .B2(KEYINPUT56), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n834_), .B1(new_n838_), .B2(new_n281_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n826_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n864_), .A2(new_n866_), .A3(new_n282_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n661_), .B1(new_n867_), .B2(new_n833_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n846_), .B1(new_n868_), .B2(KEYINPUT57), .ZN(new_n869_));
  INV_X1    g668(.A(new_n847_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n863_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT117), .B1(new_n868_), .B2(KEYINPUT57), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n849_), .A2(new_n873_), .A3(new_n850_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n862_), .B1(new_n871_), .B2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n805_), .B1(new_n876_), .B2(new_n859_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n614_), .B(new_n861_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n672_), .A2(G113gat), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n879_), .A2(G113gat), .B1(new_n877_), .B2(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT119), .ZN(G1340gat));
  INV_X1    g681(.A(new_n877_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n852_), .A2(new_n860_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n883_), .A2(KEYINPUT59), .B1(new_n884_), .B2(new_n806_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n287_), .A2(G120gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n877_), .B1(KEYINPUT60), .B2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n885_), .A2(new_n288_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(KEYINPUT60), .B2(new_n887_), .ZN(G1341gat));
  AOI21_X1  g689(.A(G127gat), .B1(new_n877_), .B2(new_n636_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n632_), .A2(G127gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n885_), .B2(new_n892_), .ZN(G1342gat));
  AOI21_X1  g692(.A(G134gat), .B1(new_n877_), .B2(new_n661_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n666_), .A2(G134gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT120), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n885_), .B2(new_n896_), .ZN(G1343gat));
  XNOR2_X1  g696(.A(KEYINPUT122), .B(G141gat), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n532_), .B1(new_n876_), .B2(new_n859_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n899_), .A2(new_n685_), .A3(new_n535_), .A4(new_n669_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT121), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n873_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n902_));
  AOI211_X1 g701(.A(KEYINPUT117), .B(KEYINPUT57), .C1(new_n843_), .C2(new_n675_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n632_), .B1(new_n904_), .B2(new_n848_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n537_), .B(new_n535_), .C1(new_n905_), .C2(new_n860_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n685_), .A4(new_n669_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n901_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n898_), .B1(new_n910_), .B2(new_n611_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n898_), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n672_), .B(new_n912_), .C1(new_n901_), .C2(new_n909_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1344gat));
  NOR2_X1   g713(.A1(new_n906_), .A2(new_n682_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n908_), .B1(new_n915_), .B2(new_n669_), .ZN(new_n916_));
  NOR4_X1   g715(.A1(new_n906_), .A2(KEYINPUT121), .A3(new_n682_), .A4(new_n668_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n288_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT123), .B(G148gat), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n910_), .A2(new_n288_), .A3(new_n919_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1345gat));
  XNOR2_X1  g722(.A(KEYINPUT61), .B(G155gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n910_), .B2(new_n636_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n924_), .ZN(new_n926_));
  AOI211_X1 g725(.A(new_n637_), .B(new_n926_), .C1(new_n901_), .C2(new_n909_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1346gat));
  AOI21_X1  g727(.A(G162gat), .B1(new_n910_), .B2(new_n661_), .ZN(new_n929_));
  INV_X1    g728(.A(G162gat), .ZN(new_n930_));
  AOI211_X1 g729(.A(new_n930_), .B(new_n724_), .C1(new_n901_), .C2(new_n909_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1347gat));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933_));
  NOR4_X1   g732(.A1(new_n669_), .A2(new_n685_), .A3(new_n537_), .A4(new_n535_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n884_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n611_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n933_), .B1(new_n937_), .B2(G169gat), .ZN(new_n938_));
  AOI211_X1 g737(.A(KEYINPUT62), .B(new_n316_), .C1(new_n936_), .C2(new_n611_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n611_), .A2(new_n319_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT124), .ZN(new_n941_));
  OAI22_X1  g740(.A1(new_n938_), .A2(new_n939_), .B1(new_n935_), .B2(new_n941_), .ZN(G1348gat));
  AOI21_X1  g741(.A(G176gat), .B1(new_n936_), .B2(new_n288_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n876_), .A2(new_n859_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n944_), .A2(new_n934_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n287_), .A2(new_n317_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n943_), .B1(new_n945_), .B2(new_n946_), .ZN(G1349gat));
  AOI21_X1  g746(.A(new_n360_), .B1(new_n945_), .B2(new_n636_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n632_), .A2(new_n353_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n936_), .B2(new_n949_), .ZN(G1350gat));
  OR3_X1    g749(.A1(new_n935_), .A2(new_n352_), .A3(new_n675_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n936_), .A2(new_n666_), .ZN(new_n952_));
  AND3_X1   g751(.A1(new_n952_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n953_));
  AOI21_X1  g752(.A(KEYINPUT125), .B1(new_n952_), .B2(G190gat), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n951_), .B1(new_n953_), .B2(new_n954_), .ZN(G1351gat));
  NOR3_X1   g754(.A1(new_n906_), .A2(new_n541_), .A3(new_n685_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n611_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g757(.A1(new_n956_), .A2(new_n288_), .ZN(new_n959_));
  XOR2_X1   g758(.A(KEYINPUT126), .B(G204gat), .Z(new_n960_));
  XNOR2_X1  g759(.A(new_n959_), .B(new_n960_), .ZN(G1353gat));
  AOI211_X1 g760(.A(KEYINPUT63), .B(G211gat), .C1(new_n956_), .C2(new_n632_), .ZN(new_n962_));
  XOR2_X1   g761(.A(KEYINPUT63), .B(G211gat), .Z(new_n963_));
  AND3_X1   g762(.A1(new_n956_), .A2(new_n632_), .A3(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n962_), .A2(new_n964_), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n956_), .B2(new_n661_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n666_), .A2(G218gat), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(KEYINPUT127), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n966_), .B1(new_n956_), .B2(new_n968_), .ZN(G1355gat));
endmodule


