//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n962_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n969_, new_n970_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_;
  XNOR2_X1  g000(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT95), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT25), .B(G183gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT23), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n207_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n208_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT92), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n209_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n216_), .A2(new_n217_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n213_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n212_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n214_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT93), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n227_), .A2(new_n229_), .A3(KEYINPUT93), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n224_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT94), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AOI211_X1 g035(.A(KEYINPUT94), .B(new_n224_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n222_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G197gat), .A2(G204gat), .ZN(new_n239_));
  OR2_X1    g038(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n239_), .B1(new_n242_), .B2(G197gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT21), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G211gat), .B(G218gat), .ZN(new_n246_));
  OR3_X1    g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n248_));
  AOI21_X1  g047(.A(G197gat), .B1(new_n240_), .B2(new_n241_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT88), .ZN(new_n250_));
  INV_X1    g049(.A(G197gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(G204gat), .ZN(new_n252_));
  INV_X1    g051(.A(G204gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n248_), .B1(new_n256_), .B2(KEYINPUT21), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n248_), .B(KEYINPUT21), .C1(new_n249_), .C2(new_n255_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n258_), .B(new_n246_), .C1(KEYINPUT21), .C2(new_n243_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n247_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n204_), .B1(new_n238_), .B2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n234_), .B(new_n235_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n258_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n246_), .B1(new_n243_), .B2(KEYINPUT21), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n256_), .A2(KEYINPUT21), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT90), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n263_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n262_), .A2(KEYINPUT95), .A3(new_n269_), .A4(new_n222_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n261_), .A2(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n225_), .A2(new_n226_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n272_), .A2(KEYINPUT82), .ZN(new_n273_));
  INV_X1    g072(.A(new_n224_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(KEYINPUT82), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n229_), .A4(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n229_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT81), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT26), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n280_), .A2(KEYINPUT79), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(KEYINPUT79), .ZN(new_n282_));
  OAI21_X1  g081(.A(G190gat), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  OR3_X1    g082(.A1(new_n280_), .A2(KEYINPUT78), .A3(G190gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT78), .B1(new_n280_), .B2(G190gat), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n283_), .A2(new_n205_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n287_), .A2(new_n212_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n229_), .A2(KEYINPUT81), .A3(KEYINPUT24), .A4(new_n219_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n279_), .A2(new_n286_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n276_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n260_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT19), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n292_), .A2(KEYINPUT20), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n271_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G8gat), .B(G36gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G64gat), .B(G92gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n238_), .A2(new_n260_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT20), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n276_), .A2(new_n290_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(new_n269_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n295_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n298_), .A2(new_n304_), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n296_), .B1(new_n261_), .B2(new_n270_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n303_), .B1(new_n312_), .B2(new_n309_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n203_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n305_), .A2(new_n295_), .A3(new_n308_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT98), .ZN(new_n316_));
  INV_X1    g115(.A(new_n233_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT93), .B1(new_n227_), .B2(new_n229_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n274_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n222_), .A2(new_n319_), .ZN(new_n320_));
  OAI211_X1 g119(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n260_), .C2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n292_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n266_), .A2(new_n268_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(new_n247_), .A3(new_n222_), .A4(new_n319_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT97), .B1(new_n324_), .B2(KEYINPUT20), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n294_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT98), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n305_), .A2(new_n308_), .A3(new_n327_), .A4(new_n295_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n316_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT99), .B1(new_n329_), .B2(new_n303_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n311_), .A2(KEYINPUT27), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(KEYINPUT99), .A3(new_n303_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n314_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G15gat), .B(G43gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT84), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n307_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n291_), .A2(new_n337_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n335_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(G71gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n342_), .A2(new_n343_), .A3(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n339_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n346_), .B1(new_n349_), .B2(new_n341_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G113gat), .B(G120gat), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n353_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(KEYINPUT85), .A3(new_n355_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n360_), .B(KEYINPUT31), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G99gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n351_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n348_), .A2(new_n350_), .A3(new_n362_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT3), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT2), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n372_), .B1(KEYINPUT1), .B2(new_n373_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT87), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n373_), .A2(new_n377_), .A3(KEYINPUT1), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n373_), .B2(KEYINPUT1), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n367_), .B(KEYINPUT86), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n369_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n375_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT29), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n384_), .A2(KEYINPUT28), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(KEYINPUT28), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n383_), .A2(KEYINPUT29), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n260_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n387_), .A2(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(G78gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G106gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G22gat), .B(G50gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n391_), .A2(new_n392_), .A3(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n385_), .A2(new_n386_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n389_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n399_), .B1(new_n404_), .B2(new_n390_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n383_), .A2(new_n359_), .A3(new_n358_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n380_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n381_), .A2(new_n369_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n413_), .A2(new_n414_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n356_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n410_), .B1(new_n409_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n408_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n409_), .A2(new_n407_), .A3(new_n416_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G85gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT0), .B(G57gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n418_), .A2(new_n419_), .A3(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n366_), .A2(new_n406_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n334_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n405_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n404_), .A2(new_n390_), .A3(new_n399_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n304_), .A2(KEYINPUT32), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n329_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n425_), .A2(new_n427_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n298_), .A2(new_n434_), .A3(new_n310_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n427_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n409_), .A2(new_n416_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n424_), .B1(new_n442_), .B2(new_n407_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(KEYINPUT4), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n411_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n443_), .B1(new_n445_), .B2(new_n407_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n427_), .B2(new_n440_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n441_), .A2(new_n447_), .A3(new_n311_), .A4(new_n313_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n433_), .B1(new_n439_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n428_), .B1(new_n401_), .B2(new_n405_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n334_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n430_), .B1(new_n452_), .B2(new_n366_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT72), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G232gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n454_), .B1(new_n457_), .B2(KEYINPUT35), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n459_));
  INV_X1    g258(.A(G99gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n396_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT7), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT7), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n459_), .A2(new_n468_), .A3(new_n460_), .A4(new_n396_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n471_));
  OR2_X1    g270(.A1(G85gat), .A2(G92gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n470_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n471_), .B1(new_n470_), .B2(new_n474_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n470_), .A2(new_n474_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(KEYINPUT67), .A3(new_n477_), .ZN(new_n480_));
  INV_X1    g279(.A(G92gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(KEYINPUT9), .ZN(new_n482_));
  AND2_X1   g281(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n482_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n396_), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n472_), .A2(KEYINPUT9), .A3(new_n473_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n485_), .A2(new_n488_), .A3(new_n489_), .A4(new_n467_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n480_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT68), .B1(new_n478_), .B2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G29gat), .B(G36gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(KEYINPUT71), .ZN(new_n496_));
  INV_X1    g295(.A(G36gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G29gat), .ZN(new_n498_));
  INV_X1    g297(.A(G29gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G36gat), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n498_), .A2(new_n500_), .A3(KEYINPUT71), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n494_), .B1(new_n496_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n500_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(KEYINPUT71), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n493_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n479_), .A2(KEYINPUT67), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n470_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(KEYINPUT8), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT68), .ZN(new_n513_));
  INV_X1    g312(.A(new_n490_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n492_), .A2(new_n509_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n515_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n508_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n502_), .A2(KEYINPUT15), .A3(new_n507_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT35), .ZN(new_n523_));
  INV_X1    g322(.A(new_n457_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n518_), .A2(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n458_), .B1(new_n517_), .B2(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n524_), .A2(KEYINPUT72), .A3(new_n523_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n528_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G190gat), .B(G218gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT36), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n529_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n535_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT36), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT102), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G230gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT64), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n513_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n552_));
  XOR2_X1   g351(.A(G71gat), .B(G78gat), .Z(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n552_), .A2(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n548_), .A2(new_n549_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n556_), .B1(new_n492_), .B2(new_n516_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n547_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT5), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT69), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n554_), .A2(new_n567_), .A3(new_n555_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n566_), .B1(new_n571_), .B2(new_n518_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n559_), .B2(new_n566_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n492_), .A2(new_n516_), .A3(new_n556_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n546_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n560_), .B(new_n565_), .C1(new_n573_), .C2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n575_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n566_), .B(new_n557_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n572_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n565_), .B1(new_n582_), .B2(new_n560_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT13), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT13), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n577_), .B2(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G15gat), .B(G22gat), .ZN(new_n589_));
  INV_X1    g388(.A(G1gat), .ZN(new_n590_));
  INV_X1    g389(.A(G8gat), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT14), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G1gat), .B(G8gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n521_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT15), .B1(new_n502_), .B2(new_n507_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT77), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT77), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n522_), .A2(new_n600_), .A3(new_n595_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n595_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n509_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n508_), .A2(new_n595_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n604_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n605_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G169gat), .B(G197gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n606_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n612_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n595_), .B(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n624_), .A2(new_n557_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n557_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT69), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n567_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT75), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT16), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT17), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT76), .Z(new_n636_));
  NOR2_X1   g435(.A1(new_n630_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n628_), .A2(KEYINPUT75), .A3(new_n629_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n634_), .A2(KEYINPUT17), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n627_), .A2(new_n635_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n588_), .A2(new_n622_), .A3(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n453_), .A2(new_n544_), .A3(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n428_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n329_), .A2(new_n303_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n311_), .A2(KEYINPUT27), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n333_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n314_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n451_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n439_), .A2(new_n448_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n406_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n366_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n334_), .A2(new_n429_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n622_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT37), .B1(new_n538_), .B2(new_n542_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n542_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT37), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n537_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n642_), .B1(new_n659_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n588_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n658_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n665_), .A2(G1gat), .A3(new_n428_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT38), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n667_), .A2(KEYINPUT101), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n666_), .B2(KEYINPUT38), .ZN(new_n671_));
  OAI221_X1 g470(.A(new_n645_), .B1(KEYINPUT38), .B2(new_n666_), .C1(new_n669_), .C2(new_n671_), .ZN(G1324gat));
  OR3_X1    g471(.A1(new_n665_), .A2(G8gat), .A3(new_n334_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n644_), .A2(new_n334_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n591_), .B1(new_n675_), .B2(KEYINPUT103), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(new_n644_), .B2(new_n334_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n544_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n657_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n650_), .A2(new_n651_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n681_), .A2(KEYINPUT103), .A3(new_n682_), .A4(new_n643_), .ZN(new_n683_));
  AND4_X1   g482(.A1(new_n674_), .A2(new_n678_), .A3(new_n683_), .A4(G8gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n673_), .B1(new_n679_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n673_), .B(KEYINPUT40), .C1(new_n679_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1325gat));
  INV_X1    g488(.A(new_n366_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G15gat), .B1(new_n644_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT41), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n665_), .A2(G15gat), .A3(new_n690_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1326gat));
  OAI21_X1  g493(.A(G22gat), .B1(new_n644_), .B2(new_n406_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n406_), .A2(G22gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n665_), .B2(new_n698_), .ZN(G1327gat));
  INV_X1    g498(.A(new_n642_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n543_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n588_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(new_n621_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n437_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n588_), .A2(new_n700_), .A3(new_n622_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n659_), .A2(new_n662_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n453_), .B2(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n707_), .B(new_n708_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n706_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n708_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n657_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n710_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(KEYINPUT44), .A3(new_n706_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n714_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n428_), .A2(new_n499_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n705_), .B1(new_n719_), .B2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(KEYINPUT106), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n714_), .A2(new_n682_), .A3(new_n718_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G36gat), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n682_), .A2(KEYINPUT105), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n334_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n497_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n704_), .A2(new_n727_), .A3(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT45), .B1(new_n703_), .B2(new_n732_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n722_), .A2(KEYINPUT106), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n724_), .B1(new_n726_), .B2(new_n739_), .ZN(new_n740_));
  AOI211_X1 g539(.A(new_n723_), .B(new_n738_), .C1(new_n725_), .C2(G36gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1329gat));
  NAND4_X1  g541(.A1(new_n714_), .A2(new_n718_), .A3(G43gat), .A4(new_n366_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G43gat), .B1(new_n704_), .B2(new_n366_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT47), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n743_), .A2(new_n748_), .A3(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1330gat));
  AOI21_X1  g549(.A(G50gat), .B1(new_n704_), .B2(new_n433_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n433_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n719_), .B2(new_n752_), .ZN(G1331gat));
  NOR2_X1   g552(.A1(new_n657_), .A2(new_n621_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n663_), .A3(new_n588_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(G57gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n437_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n664_), .A2(new_n621_), .A3(new_n642_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n681_), .A2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT107), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(new_n437_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n762_), .B2(new_n757_), .ZN(G1332gat));
  INV_X1    g562(.A(G64gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n756_), .A2(new_n764_), .A3(new_n731_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT48), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n731_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G64gat), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT48), .B(new_n764_), .C1(new_n761_), .C2(new_n731_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(G1333gat));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n761_), .A2(new_n366_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(G71gat), .ZN(new_n773_));
  AOI211_X1 g572(.A(KEYINPUT49), .B(new_n345_), .C1(new_n761_), .C2(new_n366_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n366_), .A2(new_n345_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT108), .Z(new_n776_));
  OAI22_X1  g575(.A1(new_n773_), .A2(new_n774_), .B1(new_n755_), .B2(new_n776_), .ZN(G1334gat));
  NAND3_X1  g576(.A1(new_n756_), .A2(new_n394_), .A3(new_n433_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n761_), .A2(new_n433_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(G78gat), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT50), .B(new_n394_), .C1(new_n761_), .C2(new_n433_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(G1335gat));
  NOR3_X1   g582(.A1(new_n664_), .A2(new_n701_), .A3(new_n700_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n754_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n437_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n716_), .A2(KEYINPUT109), .A3(new_n710_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n664_), .A2(new_n621_), .A3(new_n700_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n717_), .A2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n483_), .A2(new_n484_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n428_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n787_), .B1(new_n793_), .B2(new_n795_), .ZN(G1336gat));
  NAND3_X1  g595(.A1(new_n786_), .A2(new_n481_), .A3(new_n682_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n793_), .A2(new_n731_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n481_), .ZN(G1337gat));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT51), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n366_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n785_), .B2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n792_), .A2(new_n366_), .A3(new_n789_), .A4(new_n788_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(G99gat), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n800_), .A2(KEYINPUT51), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1338gat));
  NAND3_X1  g606(.A1(new_n786_), .A2(new_n396_), .A3(new_n433_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n789_), .A2(new_n433_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n717_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n811_), .B2(G106gat), .ZN(new_n812_));
  AOI211_X1 g611(.A(KEYINPUT52), .B(new_n396_), .C1(new_n717_), .C2(new_n810_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n808_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT53), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n808_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1339gat));
  NOR3_X1   g617(.A1(new_n682_), .A2(new_n428_), .A3(new_n690_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n576_), .A2(KEYINPUT113), .A3(new_n621_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT113), .B1(new_n576_), .B2(new_n621_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n547_), .B1(new_n573_), .B2(new_n558_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n578_), .A2(new_n581_), .A3(KEYINPUT55), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n827_), .A2(KEYINPUT56), .A3(new_n564_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n827_), .B2(new_n564_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n822_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n602_), .A2(new_n604_), .A3(new_n611_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n615_), .B1(new_n610_), .B2(new_n605_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n616_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n584_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n830_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT57), .B1(new_n837_), .B2(new_n701_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  AOI211_X1 g638(.A(new_n839_), .B(new_n543_), .C1(new_n830_), .C2(new_n836_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n834_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n576_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n827_), .A2(new_n564_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n827_), .A2(KEYINPUT56), .A3(new_n564_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n843_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT58), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n843_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(KEYINPUT114), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(new_n708_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n700_), .B1(new_n841_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n664_), .A2(new_n663_), .A3(new_n622_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT112), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n664_), .A2(new_n663_), .A3(new_n622_), .A4(new_n859_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n406_), .B(new_n819_), .C1(new_n856_), .C2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G113gat), .B1(new_n865_), .B2(new_n621_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n846_), .A2(new_n847_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n835_), .B1(new_n869_), .B2(new_n822_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n839_), .B1(new_n870_), .B2(new_n543_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n837_), .A2(KEYINPUT57), .A3(new_n701_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n855_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n642_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n863_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n433_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(KEYINPUT59), .A3(new_n819_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n868_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n621_), .A2(G113gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT115), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n866_), .B1(new_n878_), .B2(new_n880_), .ZN(G1340gat));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n882_));
  AOI21_X1  g681(.A(G120gat), .B1(new_n588_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT116), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n882_), .B2(G120gat), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n865_), .B(new_n884_), .C1(new_n883_), .C2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n664_), .B1(new_n868_), .B2(new_n877_), .ZN(new_n888_));
  INV_X1    g687(.A(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(G1341gat));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n642_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n868_), .B2(new_n877_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G127gat), .B1(new_n865_), .B2(new_n700_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT117), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT59), .B1(new_n876_), .B2(new_n819_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n863_), .B1(new_n873_), .B2(new_n642_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n819_), .ZN(new_n899_));
  NOR4_X1   g698(.A1(new_n898_), .A2(new_n867_), .A3(new_n433_), .A4(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n892_), .B1(new_n897_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n891_), .B1(new_n864_), .B2(new_n642_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n896_), .A2(new_n904_), .ZN(G1342gat));
  INV_X1    g704(.A(G134gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n864_), .B2(new_n544_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT118), .B(new_n906_), .C1(new_n864_), .C2(new_n544_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n715_), .A2(new_n906_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n909_), .A2(new_n910_), .B1(new_n878_), .B2(new_n911_), .ZN(G1343gat));
  NAND2_X1  g711(.A1(new_n874_), .A2(new_n875_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n731_), .A2(new_n428_), .A3(new_n406_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n913_), .A2(new_n690_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n621_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n588_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g718(.A(KEYINPUT61), .B(G155gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT120), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT119), .B1(new_n915_), .B2(new_n700_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n913_), .A2(new_n690_), .A3(new_n914_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n924_), .A2(new_n925_), .A3(new_n642_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n922_), .B1(new_n923_), .B2(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n915_), .A2(KEYINPUT119), .A3(new_n700_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n925_), .B1(new_n924_), .B2(new_n642_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n928_), .A2(new_n929_), .A3(new_n921_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n927_), .A2(new_n930_), .ZN(G1346gat));
  OR3_X1    g730(.A1(new_n924_), .A2(G162gat), .A3(new_n544_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G162gat), .B1(new_n924_), .B2(new_n715_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1347gat));
  NAND3_X1  g733(.A1(new_n731_), .A2(new_n428_), .A3(new_n366_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n935_), .A2(KEYINPUT121), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(KEYINPUT121), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n939_), .A2(new_n621_), .A3(new_n876_), .ZN(new_n940_));
  XOR2_X1   g739(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n941_));
  AND3_X1   g740(.A1(new_n940_), .A2(G169gat), .A3(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(G169gat), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n939_), .A2(new_n876_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n621_), .A2(new_n225_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(KEYINPUT123), .ZN(new_n946_));
  OAI22_X1  g745(.A1(new_n942_), .A2(new_n943_), .B1(new_n944_), .B2(new_n946_), .ZN(G1348gat));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n948_), .B1(new_n898_), .B2(new_n433_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n949_), .A2(new_n939_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n876_), .A2(KEYINPUT125), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n664_), .A2(new_n226_), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .A4(new_n953_), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n952_), .A2(new_n949_), .A3(new_n939_), .A4(new_n953_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(KEYINPUT126), .ZN(new_n956_));
  NOR4_X1   g755(.A1(new_n938_), .A2(new_n898_), .A3(new_n433_), .A4(new_n664_), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT124), .B1(new_n957_), .B2(G176gat), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n959_), .B(new_n226_), .C1(new_n944_), .C2(new_n664_), .ZN(new_n960_));
  AOI22_X1  g759(.A1(new_n954_), .A2(new_n956_), .B1(new_n958_), .B2(new_n960_), .ZN(G1349gat));
  NOR3_X1   g760(.A1(new_n944_), .A2(new_n205_), .A3(new_n642_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n950_), .A2(new_n700_), .A3(new_n952_), .ZN(new_n963_));
  INV_X1    g762(.A(G183gat), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n962_), .B1(new_n963_), .B2(new_n964_), .ZN(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n944_), .B2(new_n715_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n680_), .A2(new_n206_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n944_), .B2(new_n967_), .ZN(G1351gat));
  NOR2_X1   g767(.A1(new_n898_), .A2(new_n366_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n450_), .B1(new_n728_), .B2(new_n730_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n971_), .A2(new_n622_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(new_n251_), .ZN(G1352gat));
  INV_X1    g772(.A(new_n971_), .ZN(new_n974_));
  AOI21_X1  g773(.A(G204gat), .B1(new_n974_), .B2(new_n588_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n971_), .A2(new_n664_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n975_), .B1(new_n242_), .B2(new_n976_), .ZN(G1353gat));
  AOI21_X1  g776(.A(new_n642_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(KEYINPUT127), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n971_), .A2(new_n979_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n980_), .B(new_n981_), .ZN(G1354gat));
  OR3_X1    g781(.A1(new_n971_), .A2(G218gat), .A3(new_n544_), .ZN(new_n983_));
  OAI21_X1  g782(.A(G218gat), .B1(new_n971_), .B2(new_n715_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n983_), .A2(new_n984_), .ZN(G1355gat));
endmodule


