//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_;
  NAND3_X1  g000(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT83), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT83), .ZN(new_n204_));
  NAND4_X1  g003(.A1(new_n204_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G141gat), .ZN(new_n209_));
  INV_X1    g008(.A(G148gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT3), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(G141gat), .B2(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n206_), .A2(new_n208_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT84), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n207_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT84), .A3(new_n206_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n217_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n220_), .A2(KEYINPUT1), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n209_), .A2(new_n210_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n218_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G127gat), .B(G134gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G113gat), .ZN(new_n231_));
  INV_X1    g030(.A(G120gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G225gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n229_), .B(new_n233_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n235_), .B(new_n237_), .C1(new_n238_), .C2(new_n234_), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n229_), .B(new_n233_), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n236_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT0), .B(G57gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G85gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(G1gat), .B(G29gat), .Z(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  NOR2_X1   g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n246_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G85gat), .B(G92gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT65), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G99gat), .A2(G106gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT6), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n255_));
  OR3_X1    g054(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT8), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT9), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n251_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G92gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(KEYINPUT9), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n264_), .A2(G92gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(G85gat), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT10), .B(G99gat), .Z(new_n269_));
  INV_X1    g068(.A(G106gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n263_), .A2(new_n268_), .A3(new_n254_), .A4(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n252_), .A2(KEYINPUT66), .A3(new_n257_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT8), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT66), .B1(new_n252_), .B2(new_n257_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n261_), .B(new_n272_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G57gat), .B(G64gat), .Z(new_n279_));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G57gat), .B(G64gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT11), .ZN(new_n283_));
  XOR2_X1   g082(.A(G71gat), .B(G78gat), .Z(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n283_), .A2(new_n284_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT68), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n258_), .A2(new_n259_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(KEYINPUT8), .A3(new_n273_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n291_), .A2(KEYINPUT67), .A3(new_n261_), .A4(new_n272_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n278_), .A2(new_n289_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n285_), .A2(new_n286_), .A3(KEYINPUT69), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT69), .B1(new_n285_), .B2(new_n286_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n276_), .A2(KEYINPUT12), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n276_), .A2(new_n298_), .A3(KEYINPUT70), .A4(KEYINPUT12), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G230gat), .A2(G233gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n278_), .A2(new_n292_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n288_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n295_), .A2(new_n303_), .A3(new_n304_), .A4(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n293_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n289_), .B1(new_n278_), .B2(new_n292_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G120gat), .B(G148gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT72), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G176gat), .B(G204gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n307_), .A2(new_n311_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n307_), .B2(new_n311_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT13), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G1gat), .A2(G8gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT14), .ZN(new_n324_));
  INV_X1    g123(.A(G15gat), .ZN(new_n325_));
  INV_X1    g124(.A(G22gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G15gat), .A2(G22gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n324_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT74), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n331_), .B(new_n324_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G1gat), .B(G8gat), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n330_), .A2(new_n334_), .A3(new_n332_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G29gat), .B(G36gat), .ZN(new_n339_));
  INV_X1    g138(.A(G43gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G50gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n339_), .B(G43gat), .ZN(new_n343_));
  INV_X1    g142(.A(G50gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n338_), .A2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n336_), .A2(new_n342_), .A3(new_n345_), .A4(new_n337_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(KEYINPUT76), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G229gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n338_), .A2(new_n346_), .A3(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n342_), .A2(new_n345_), .A3(KEYINPUT15), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT15), .B1(new_n342_), .B2(new_n345_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n338_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n350_), .A3(new_n348_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT77), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G113gat), .B(G141gat), .ZN(new_n360_));
  INV_X1    g159(.A(G169gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G197gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n359_), .B(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT13), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n322_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G8gat), .B(G36gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT19), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n378_), .A2(new_n379_), .A3(G197gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(new_n363_), .B2(G204gat), .ZN(new_n382_));
  INV_X1    g181(.A(G204gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT21), .B1(new_n380_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G211gat), .B(G218gat), .Z(new_n389_));
  NOR2_X1   g188(.A1(new_n383_), .A2(G197gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT88), .B(G204gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(G197gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT21), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n389_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT89), .B(KEYINPUT21), .C1(new_n380_), .C2(new_n385_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n388_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n393_), .B1(new_n389_), .B2(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n391_), .A2(G197gat), .ZN(new_n399_));
  OAI221_X1 g198(.A(new_n398_), .B1(new_n397_), .B2(new_n389_), .C1(new_n399_), .C2(new_n390_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G176gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n361_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G169gat), .A2(G176gat), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n403_), .A2(KEYINPUT24), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT23), .ZN(new_n406_));
  INV_X1    g205(.A(G183gat), .ZN(new_n407_));
  INV_X1    g206(.A(G190gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n403_), .A2(KEYINPUT24), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n405_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(G190gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT25), .B(G183gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G190gat), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n416_), .B(new_n417_), .C1(new_n418_), .C2(new_n414_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n407_), .A2(new_n408_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n409_), .A2(new_n421_), .A3(new_n410_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT79), .ZN(new_n423_));
  INV_X1    g222(.A(new_n404_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT22), .B(G169gat), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n425_), .B2(new_n402_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n409_), .A2(new_n421_), .A3(new_n427_), .A4(new_n410_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n420_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT80), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT80), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n420_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n401_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n418_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n417_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n413_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n426_), .A2(new_n422_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT99), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n401_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n377_), .B1(new_n436_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n401_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n440_), .A2(KEYINPUT95), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n440_), .A2(KEYINPUT95), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n439_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n396_), .A2(new_n400_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n435_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n445_), .A2(new_n377_), .A3(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n374_), .B1(new_n444_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n377_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n431_), .A2(new_n433_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n449_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n448_), .A2(new_n449_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT20), .A4(new_n377_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n458_), .A3(new_n373_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n452_), .A2(KEYINPUT27), .A3(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n377_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n434_), .A2(new_n461_), .A3(new_n435_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n374_), .B1(new_n462_), .B2(new_n453_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT27), .B1(new_n463_), .B2(new_n459_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT100), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n464_), .A2(new_n465_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n250_), .B(new_n460_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n455_), .A2(new_n233_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n455_), .A2(new_n233_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT31), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G227gat), .A2(G233gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n471_), .A2(new_n472_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G71gat), .B(G99gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT30), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G15gat), .B(G43gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OR3_X1    g283(.A1(new_n478_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G78gat), .B(G106gat), .Z(new_n489_));
  AND3_X1   g288(.A1(new_n222_), .A2(KEYINPUT84), .A3(new_n206_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT84), .B1(new_n222_), .B2(new_n206_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n220_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT29), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n449_), .B1(new_n494_), .B2(KEYINPUT86), .ZN(new_n495_));
  INV_X1    g294(.A(G228gat), .ZN(new_n496_));
  INV_X1    g295(.A(G233gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT29), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n500_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n499_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n495_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n494_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(KEYINPUT91), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n449_), .A3(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n509_), .A2(KEYINPUT92), .A3(new_n498_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT92), .B1(new_n509_), .B2(new_n498_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n489_), .B(new_n505_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n224_), .A2(new_n500_), .A3(new_n228_), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n514_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G22gat), .B(G50gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n515_), .A2(new_n518_), .A3(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n522_), .A2(KEYINPUT93), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n512_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT91), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n526_));
  AOI211_X1 g325(.A(new_n506_), .B(new_n500_), .C1(new_n224_), .C2(new_n228_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n401_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n525_), .B1(new_n528_), .B2(new_n499_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n509_), .A2(KEYINPUT92), .A3(new_n498_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n489_), .B1(new_n531_), .B2(new_n505_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n489_), .ZN(new_n533_));
  AOI211_X1 g332(.A(new_n533_), .B(new_n504_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n524_), .B1(new_n535_), .B2(new_n523_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n522_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n504_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n538_), .A2(KEYINPUT94), .A3(new_n489_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n505_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n540_), .B1(new_n541_), .B2(new_n533_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n537_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n488_), .B1(new_n536_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n533_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n523_), .A3(new_n512_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n512_), .A2(new_n523_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT94), .B1(new_n538_), .B2(new_n489_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n540_), .A3(new_n533_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n522_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n548_), .A2(new_n551_), .A3(new_n487_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n470_), .B1(new_n544_), .B2(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(KEYINPUT32), .B(new_n373_), .C1(new_n444_), .C2(new_n451_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n373_), .A2(KEYINPUT32), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n454_), .A2(new_n458_), .A3(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n554_), .B(new_n556_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n462_), .A2(new_n453_), .A3(new_n374_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n373_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT97), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n463_), .A2(new_n459_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n242_), .B2(new_n246_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n239_), .A2(new_n241_), .A3(new_n248_), .A4(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n240_), .A2(new_n237_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n235_), .B1(new_n238_), .B2(new_n234_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n246_), .B(new_n568_), .C1(new_n569_), .C2(new_n237_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n565_), .A2(new_n567_), .A3(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n557_), .B1(new_n563_), .B2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n572_), .B(new_n488_), .C1(new_n551_), .C2(new_n548_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n368_), .B1(new_n553_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n346_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n355_), .A2(new_n356_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n305_), .A2(new_n575_), .B1(new_n576_), .B2(new_n276_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(KEYINPUT35), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n579_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT35), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n577_), .B2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(G134gat), .ZN(new_n588_));
  INV_X1    g387(.A(G162gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT36), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n581_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n581_), .B2(new_n586_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT73), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(KEYINPUT73), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n593_), .A2(new_n596_), .A3(KEYINPUT73), .A4(new_n598_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n338_), .B(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(new_n298_), .Z(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT16), .B(G183gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(G211gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n606_), .B(new_n288_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n613_), .B(KEYINPUT17), .Z(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n604_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n574_), .A2(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT101), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT101), .ZN(new_n622_));
  AOI211_X1 g421(.A(G1gat), .B(new_n250_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT38), .Z(new_n624_));
  INV_X1    g423(.A(new_n618_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n597_), .B(KEYINPUT102), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n574_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G1gat), .B1(new_n627_), .B2(new_n250_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(G1324gat));
  INV_X1    g428(.A(new_n468_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n466_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n460_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n627_), .A2(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(G8gat), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n634_), .B2(G8gat), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(G8gat), .B1(new_n621_), .B2(new_n622_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n639_), .A2(new_n640_), .A3(new_n632_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n639_), .B2(new_n632_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n638_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT105), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n638_), .B(new_n645_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n627_), .B2(new_n488_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT41), .Z(new_n651_));
  INV_X1    g450(.A(new_n620_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n325_), .A3(new_n487_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT107), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(G1326gat));
  NOR2_X1   g454(.A1(new_n548_), .A2(new_n551_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G22gat), .B1(new_n627_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT42), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n652_), .A2(new_n326_), .A3(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n553_), .A2(new_n573_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n368_), .A2(new_n625_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n597_), .A3(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n665_), .A2(G29gat), .A3(new_n250_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n663_), .B2(new_n604_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n487_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n543_), .A2(new_n488_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n469_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n573_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n604_), .B(new_n668_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT44), .B(new_n664_), .C1(new_n669_), .C2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n664_), .B1(new_n669_), .B2(new_n675_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n664_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n604_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT43), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n682_), .B1(new_n684_), .B2(new_n674_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT108), .B1(new_n685_), .B2(KEYINPUT44), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n677_), .B1(new_n681_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n250_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(G29gat), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n662_), .B(new_n667_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT109), .B1(new_n692_), .B2(new_n666_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1328gat));
  INV_X1    g493(.A(KEYINPUT111), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(KEYINPUT112), .B2(KEYINPUT46), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n633_), .B1(new_n685_), .B2(KEYINPUT44), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n679_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n685_), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G36gat), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n665_), .A2(G36gat), .A3(new_n633_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n696_), .B1(new_n701_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n676_), .A2(new_n632_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n686_), .B2(new_n681_), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT111), .B(new_n704_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT112), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n705_), .B1(new_n710_), .B2(new_n711_), .ZN(G1329gat));
  NAND2_X1  g511(.A1(KEYINPUT113), .A2(G43gat), .ZN(new_n713_));
  OR2_X1    g512(.A1(KEYINPUT113), .A2(G43gat), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n713_), .B(new_n714_), .C1(new_n665_), .C2(new_n488_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT114), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n488_), .A2(new_n340_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n687_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(G1330gat));
  AND2_X1   g519(.A1(new_n687_), .A2(new_n656_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n656_), .A2(new_n344_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT115), .Z(new_n723_));
  OAI22_X1  g522(.A1(new_n721_), .A2(new_n344_), .B1(new_n665_), .B2(new_n723_), .ZN(G1331gat));
  AOI21_X1  g523(.A(new_n365_), .B1(new_n322_), .B2(new_n367_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n663_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n619_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n688_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n250_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(G57gat), .B2(new_n731_), .ZN(G1332gat));
  OAI21_X1  g531(.A(G64gat), .B1(new_n730_), .B2(new_n633_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT48), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n633_), .A2(G64gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n727_), .B2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n730_), .B2(new_n488_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT49), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n488_), .A2(G71gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n727_), .B2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n730_), .B2(new_n657_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n727_), .A2(G78gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n657_), .B2(new_n743_), .ZN(G1335gat));
  NAND4_X1  g543(.A1(new_n663_), .A2(new_n618_), .A3(new_n597_), .A4(new_n725_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n688_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n725_), .A2(new_n618_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT116), .Z(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n669_), .B2(new_n675_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(new_n250_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n747_), .B1(new_n751_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g551(.A(G92gat), .B1(new_n746_), .B2(new_n632_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n750_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n267_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n633_), .B1(new_n755_), .B2(new_n265_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n754_), .B2(new_n756_), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n746_), .A2(new_n269_), .A3(new_n487_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT117), .ZN(new_n759_));
  INV_X1    g558(.A(G99gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n754_), .B2(new_n487_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(G1338gat));
  OAI21_X1  g563(.A(G106gat), .B1(new_n750_), .B2(new_n657_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n745_), .A2(G106gat), .A3(new_n657_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT118), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT52), .B(G106gat), .C1(new_n750_), .C2(new_n657_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g571(.A1(new_n632_), .A2(new_n250_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n365_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT119), .B1(new_n319_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT119), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n318_), .A2(new_n778_), .A3(new_n365_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n310_), .B1(new_n294_), .B2(new_n293_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n304_), .B1(new_n781_), .B2(new_n303_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n307_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n295_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(new_n783_), .A3(new_n308_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n317_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n791_), .B(new_n317_), .C1(new_n784_), .C2(new_n787_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n780_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n351_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n350_), .B1(new_n357_), .B2(new_n348_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n364_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n364_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n354_), .A2(new_n358_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n321_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n793_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n597_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n775_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n597_), .B(new_n774_), .C1(new_n793_), .C2(new_n801_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n317_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(KEYINPUT56), .ZN(new_n809_));
  AND4_X1   g608(.A1(new_n304_), .A2(new_n295_), .A3(new_n303_), .A4(new_n306_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n785_), .A2(new_n308_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(KEYINPUT55), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n789_), .B1(new_n812_), .B2(new_n786_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT121), .A3(new_n791_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n789_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n809_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n319_), .A2(new_n799_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(KEYINPUT58), .A3(new_n817_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n604_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n625_), .B1(new_n806_), .B2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n602_), .A2(new_n625_), .A3(new_n776_), .A4(new_n603_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n322_), .A2(new_n367_), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n824_), .A2(KEYINPUT54), .A3(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT54), .B1(new_n824_), .B2(new_n825_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n544_), .B(new_n773_), .C1(new_n823_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n365_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n816_), .A2(KEYINPUT58), .A3(new_n817_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT58), .B1(new_n816_), .B2(new_n817_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n604_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n777_), .A2(new_n779_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n813_), .A2(new_n791_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n815_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n803_), .B1(new_n841_), .B2(new_n800_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n774_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n802_), .A2(new_n803_), .A3(new_n775_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n618_), .B1(new_n838_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n670_), .B1(new_n846_), .B2(new_n828_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT59), .A3(new_n773_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n776_), .B1(new_n834_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n832_), .B1(new_n849_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g649(.A(new_n825_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n232_), .B1(new_n851_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT122), .B1(new_n232_), .B2(KEYINPUT60), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n830_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n852_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n851_), .B1(new_n834_), .B2(new_n848_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n232_), .ZN(G1341gat));
  AOI21_X1  g657(.A(G127gat), .B1(new_n831_), .B2(new_n625_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n618_), .B1(new_n834_), .B2(new_n848_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g660(.A(new_n626_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G134gat), .B1(new_n831_), .B2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n837_), .B1(new_n834_), .B2(new_n848_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n806_), .A2(new_n822_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n829_), .B1(new_n866_), .B2(new_n618_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n773_), .A2(new_n552_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT123), .Z(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n867_), .A2(KEYINPUT124), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n846_), .A2(new_n828_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n869_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n365_), .B1(new_n871_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G141gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT124), .B1(new_n867_), .B2(new_n870_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n873_), .A2(new_n872_), .A3(new_n869_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n209_), .A3(new_n365_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n880_), .ZN(G1344gat));
  OAI21_X1  g680(.A(new_n825_), .B1(new_n871_), .B2(new_n874_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT125), .B(G148gat), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n879_), .A2(new_n825_), .A3(new_n883_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1345gat));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n879_), .B2(new_n625_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n888_), .ZN(new_n890_));
  AOI211_X1 g689(.A(new_n618_), .B(new_n890_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n879_), .B2(new_n862_), .ZN(new_n893_));
  AOI211_X1 g692(.A(new_n589_), .B(new_n837_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n633_), .A2(new_n688_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n544_), .B(new_n896_), .C1(new_n823_), .C2(new_n829_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(KEYINPUT126), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n847_), .B2(new_n896_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n365_), .B(new_n425_), .C1(new_n898_), .C2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n847_), .A2(new_n365_), .A3(new_n896_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n902_), .A2(new_n903_), .A3(G169gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n902_), .B2(G169gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n901_), .B1(new_n904_), .B2(new_n905_), .ZN(G1348gat));
  OAI21_X1  g705(.A(G176gat), .B1(new_n897_), .B2(new_n851_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n402_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n851_), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n897_), .A2(KEYINPUT126), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n847_), .A2(new_n899_), .A3(new_n896_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n618_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n847_), .A2(new_n625_), .A3(new_n896_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n912_), .A2(new_n438_), .B1(new_n407_), .B2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(new_n862_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n837_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n916_));
  OAI22_X1  g715(.A1(new_n915_), .A2(new_n437_), .B1(new_n916_), .B2(new_n408_), .ZN(G1351gat));
  OAI211_X1 g716(.A(new_n552_), .B(new_n896_), .C1(new_n823_), .C2(new_n829_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n776_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(new_n363_), .ZN(G1352gat));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n851_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n391_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n922_), .B1(new_n383_), .B2(new_n921_), .ZN(G1353gat));
  NOR2_X1   g722(.A1(new_n918_), .A2(new_n618_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n926_));
  INV_X1    g725(.A(G211gat), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(new_n927_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n924_), .A2(new_n925_), .A3(new_n928_), .A4(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n671_), .B1(new_n846_), .B2(new_n828_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n932_), .A2(new_n625_), .A3(new_n896_), .A4(new_n928_), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT127), .B1(new_n933_), .B2(new_n929_), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n926_), .B(new_n927_), .C1(new_n918_), .C2(new_n618_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n931_), .A2(new_n934_), .A3(new_n935_), .ZN(G1354gat));
  NOR2_X1   g735(.A1(new_n918_), .A2(new_n626_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(G218gat), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n918_), .A2(new_n837_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(G218gat), .B2(new_n939_), .ZN(G1355gat));
endmodule


