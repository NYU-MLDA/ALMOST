//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G71gat), .B(G78gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  INV_X1    g004(.A(G64gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G57gat), .ZN(new_n207_));
  INV_X1    g006(.A(G57gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G64gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n209_), .A3(KEYINPUT11), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n205_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n204_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(G231gat), .A2(G233gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT78), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217_));
  INV_X1    g016(.A(G1gat), .ZN(new_n218_));
  INV_X1    g017(.A(G8gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT14), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G1gat), .B(G8gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n216_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G127gat), .B(G155gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT16), .ZN(new_n227_));
  XOR2_X1   g026(.A(G183gat), .B(G211gat), .Z(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n230_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n225_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT80), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n225_), .B(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n237_), .A2(KEYINPUT79), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n231_), .B1(new_n237_), .B2(KEYINPUT79), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n235_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G85gat), .B(G92gat), .Z(new_n242_));
  NAND2_X1  g041(.A1(G99gat), .A2(G106gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246_));
  INV_X1    g045(.A(G99gat), .ZN(new_n247_));
  INV_X1    g046(.A(G106gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n242_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT8), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT8), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n254_), .B(new_n242_), .C1(new_n245_), .C2(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257_));
  INV_X1    g056(.A(G85gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259_));
  INV_X1    g058(.A(G92gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n257_), .B1(new_n263_), .B2(KEYINPUT9), .ZN(new_n264_));
  INV_X1    g063(.A(new_n262_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(G85gat), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT9), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(KEYINPUT66), .A3(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT67), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(G85gat), .B2(G92gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n273_), .B2(new_n270_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n264_), .A2(new_n269_), .A3(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(KEYINPUT64), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n280_));
  INV_X1    g079(.A(new_n278_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(new_n281_), .B2(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n245_), .B1(new_n283_), .B2(new_n248_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n275_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G43gat), .B(G50gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G36gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G29gat), .ZN(new_n289_));
  INV_X1    g088(.A(G29gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G36gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n291_), .A3(KEYINPUT74), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT74), .B1(new_n289_), .B2(new_n291_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n287_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(new_n291_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n292_), .A3(new_n286_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n256_), .A2(new_n285_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT15), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n295_), .A2(new_n299_), .A3(KEYINPUT15), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n253_), .A2(new_n255_), .B1(new_n275_), .B2(new_n284_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n301_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n308_));
  NAND2_X1  g107(.A1(G232gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT35), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n307_), .A2(KEYINPUT75), .A3(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n310_), .B(KEYINPUT35), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n301_), .B(new_n318_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT77), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n256_), .A2(new_n285_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(new_n304_), .A3(new_n303_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n301_), .A4(new_n318_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G190gat), .B(G218gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G134gat), .B(G162gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(KEYINPUT36), .A3(new_n329_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n315_), .A2(new_n316_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n329_), .A2(KEYINPUT36), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n331_), .A2(KEYINPUT76), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n332_), .B1(new_n331_), .B2(KEYINPUT76), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n330_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT37), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT37), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n337_), .B(new_n330_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n241_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n256_), .A2(new_n285_), .A3(new_n213_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G230gat), .A2(G233gat), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n213_), .B1(new_n256_), .B2(new_n285_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n213_), .A2(KEYINPUT68), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n236_), .B(new_n204_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT12), .A3(new_n351_), .ZN(new_n352_));
  OAI22_X1  g151(.A1(new_n349_), .A2(KEYINPUT12), .B1(new_n306_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n342_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n353_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n355_), .B(KEYINPUT70), .C1(new_n347_), .C2(new_n346_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n343_), .ZN(new_n357_));
  OAI211_X1 g156(.A(G230gat), .B(G233gat), .C1(new_n357_), .C2(new_n349_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G120gat), .B(G148gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(G176gat), .B(G204gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n359_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n354_), .A2(new_n356_), .A3(new_n358_), .A4(new_n364_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT13), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n369_), .A2(KEYINPUT72), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(KEYINPUT72), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n224_), .A2(new_n300_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n223_), .A2(new_n299_), .A3(new_n295_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G229gat), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n303_), .A2(new_n223_), .A3(new_n304_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n224_), .B2(new_n300_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n375_), .A2(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G113gat), .B(G141gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G169gat), .B(G197gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  AND3_X1   g182(.A1(new_n380_), .A2(KEYINPUT82), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT82), .B1(new_n380_), .B2(new_n383_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n375_), .A2(new_n377_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n378_), .A2(new_n379_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n383_), .B1(new_n389_), .B2(KEYINPUT81), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(KEYINPUT81), .B2(new_n389_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n372_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(KEYINPUT1), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n396_), .B2(KEYINPUT1), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT90), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n398_), .B2(new_n397_), .ZN(new_n400_));
  OR2_X1    g199(.A1(G141gat), .A2(G148gat), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n401_), .A2(KEYINPUT89), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(KEYINPUT89), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n402_), .A2(new_n403_), .B1(G141gat), .B2(G148gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT91), .ZN(new_n406_));
  INV_X1    g205(.A(new_n396_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT92), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n401_), .B(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n411_), .B(KEYINPUT2), .Z(new_n412_));
  OAI211_X1 g211(.A(new_n394_), .B(new_n407_), .C1(new_n410_), .C2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G127gat), .B(G134gat), .Z(new_n415_));
  XOR2_X1   g214(.A(G113gat), .B(G120gat), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT87), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n415_), .A2(new_n416_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n414_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n417_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT102), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n406_), .A2(new_n413_), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n422_), .A2(KEYINPUT4), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n414_), .A2(new_n429_), .A3(new_n421_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n427_), .A3(new_n425_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G85gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT0), .B(G57gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n431_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n414_), .A2(KEYINPUT29), .ZN(new_n444_));
  XOR2_X1   g243(.A(G211gat), .B(G218gat), .Z(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT95), .B(G204gat), .Z(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT94), .B(G197gat), .Z(new_n447_));
  OAI22_X1  g246(.A1(G197gat), .A2(new_n446_), .B1(new_n447_), .B2(G204gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n445_), .B1(new_n448_), .B2(KEYINPUT21), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(G197gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT96), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n447_), .A2(G204gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT97), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n449_), .B1(new_n454_), .B2(KEYINPUT21), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT21), .A3(new_n445_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n444_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G233gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT93), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(G228gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(G228gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n459_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n458_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n464_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n444_), .A2(new_n457_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n443_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n465_), .A2(new_n467_), .A3(new_n443_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n414_), .A2(KEYINPUT29), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G22gat), .B(G50gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT28), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n472_), .B(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n468_), .B2(KEYINPUT98), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n469_), .A2(new_n470_), .A3(KEYINPUT98), .A4(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G183gat), .A2(G190gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n482_), .A2(KEYINPUT23), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  MUX2_X1   g284(.A(new_n483_), .B(new_n485_), .S(KEYINPUT85), .Z(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT83), .B(G183gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT25), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n489_), .B1(KEYINPUT25), .B2(G183gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT26), .B(G190gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(G169gat), .B2(G176gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  OR3_X1    g294(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n486_), .A2(new_n492_), .A3(new_n495_), .A4(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n482_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(KEYINPUT23), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(new_n498_), .B2(new_n481_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(G190gat), .B2(new_n488_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(G169gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n497_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT86), .B(G15gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n497_), .B2(new_n504_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n509_), .A2(new_n420_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G71gat), .B(G99gat), .ZN(new_n514_));
  INV_X1    g313(.A(G43gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT30), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT31), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n420_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n513_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n513_), .B2(new_n519_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n480_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(KEYINPUT88), .A3(new_n520_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n479_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n521_), .A2(new_n522_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n477_), .A2(new_n478_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n441_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT105), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n486_), .B1(G183gat), .B2(G190gat), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n532_), .A2(new_n503_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n500_), .A2(new_n496_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT100), .ZN(new_n535_));
  INV_X1    g334(.A(new_n491_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT25), .B(G183gat), .Z(new_n537_));
  OAI21_X1  g336(.A(new_n495_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n531_), .B1(new_n533_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n457_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n532_), .A2(new_n503_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n542_), .B(KEYINPUT105), .C1(new_n535_), .C2(new_n538_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n540_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n457_), .A2(new_n505_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT101), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n457_), .A2(KEYINPUT101), .A3(new_n505_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n544_), .A2(KEYINPUT20), .A3(new_n547_), .A4(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G226gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT19), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT106), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT106), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n554_), .A3(new_n551_), .ZN(new_n555_));
  OAI211_X1 g354(.A(KEYINPUT99), .B(KEYINPUT20), .C1(new_n457_), .C2(new_n505_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n457_), .B1(new_n533_), .B2(new_n539_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n551_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT20), .B1(new_n457_), .B2(new_n505_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT99), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT107), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n558_), .A2(KEYINPUT107), .A3(new_n559_), .A4(new_n562_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n553_), .A2(new_n555_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G8gat), .B(G36gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT18), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G64gat), .B(G92gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT108), .B1(new_n567_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT108), .ZN(new_n573_));
  INV_X1    g372(.A(new_n571_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n565_), .A2(new_n566_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n549_), .A2(new_n554_), .A3(new_n551_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n554_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n573_), .B(new_n574_), .C1(new_n575_), .C2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n533_), .A2(new_n539_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n551_), .B1(new_n580_), .B2(new_n541_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n581_), .A2(new_n547_), .A3(KEYINPUT20), .A4(new_n548_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n558_), .A2(new_n562_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n571_), .B(new_n582_), .C1(new_n583_), .C2(new_n559_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n584_), .A2(KEYINPUT27), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n572_), .A2(new_n579_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n559_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n582_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n574_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT27), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n530_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n526_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n479_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n440_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT104), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n426_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n422_), .A2(new_n428_), .A3(new_n425_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n438_), .A3(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n584_), .A2(new_n589_), .A3(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT33), .A4(new_n437_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT103), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n597_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n582_), .B1(new_n583_), .B2(new_n559_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n571_), .A2(KEYINPUT32), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n441_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n567_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n610_), .B2(new_n608_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n594_), .B1(new_n605_), .B2(new_n611_), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n341_), .B(new_n393_), .C1(new_n592_), .C2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n218_), .A3(new_n441_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n614_), .A2(KEYINPUT109), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(KEYINPUT109), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n615_), .A2(KEYINPUT38), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT38), .B1(new_n615_), .B2(new_n616_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n393_), .A2(new_n240_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n335_), .B1(new_n592_), .B2(new_n612_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n218_), .B1(new_n621_), .B2(new_n441_), .ZN(new_n622_));
  OR3_X1    g421(.A1(new_n617_), .A2(new_n618_), .A3(new_n622_), .ZN(G1324gat));
  NAND2_X1  g422(.A1(new_n586_), .A2(new_n591_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n613_), .A2(new_n219_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n219_), .B1(KEYINPUT110), .B2(KEYINPUT39), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT110), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n625_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(KEYINPUT40), .B(new_n625_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1325gat));
  INV_X1    g436(.A(G15gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n621_), .B2(new_n593_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT41), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n613_), .A2(new_n638_), .A3(new_n593_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n621_), .B2(new_n479_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT42), .Z(new_n645_));
  NAND3_X1  g444(.A1(new_n613_), .A2(new_n643_), .A3(new_n479_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n393_), .A2(new_n241_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n592_), .A2(new_n612_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(new_n339_), .ZN(new_n651_));
  AOI211_X1 g450(.A(KEYINPUT43), .B(new_n340_), .C1(new_n592_), .C2(new_n612_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT44), .B(new_n648_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n655_), .A2(G29gat), .A3(new_n441_), .A4(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n393_), .B1(new_n592_), .B2(new_n612_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n335_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n241_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n441_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n290_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n657_), .A2(new_n663_), .ZN(G1328gat));
  NAND3_X1  g463(.A1(new_n655_), .A2(new_n624_), .A3(new_n656_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G36gat), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n658_), .A2(new_n288_), .A3(new_n624_), .A4(new_n660_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT45), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n666_), .A2(KEYINPUT46), .A3(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1329gat));
  NAND4_X1  g472(.A1(new_n655_), .A2(G43gat), .A3(new_n528_), .A4(new_n656_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n515_), .B1(new_n661_), .B2(new_n526_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g476(.A1(new_n655_), .A2(G50gat), .A3(new_n479_), .A4(new_n656_), .ZN(new_n678_));
  INV_X1    g477(.A(G50gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n479_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n661_), .B2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n678_), .A2(new_n681_), .ZN(G1331gat));
  INV_X1    g481(.A(new_n372_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n392_), .ZN(new_n684_));
  AND4_X1   g483(.A1(new_n241_), .A2(new_n620_), .A3(new_n683_), .A4(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n208_), .B1(new_n685_), .B2(new_n441_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n392_), .B1(new_n592_), .B2(new_n612_), .ZN(new_n687_));
  AND4_X1   g486(.A1(new_n241_), .A2(new_n687_), .A3(new_n340_), .A4(new_n683_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n662_), .A2(G57gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT111), .ZN(G1332gat));
  AOI21_X1  g490(.A(new_n206_), .B1(new_n685_), .B2(new_n624_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n688_), .A2(new_n206_), .A3(new_n624_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1333gat));
  INV_X1    g495(.A(G71gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n685_), .B2(new_n593_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT49), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n688_), .A2(new_n697_), .A3(new_n593_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1334gat));
  INV_X1    g500(.A(G78gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n685_), .B2(new_n479_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT50), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n688_), .A2(new_n702_), .A3(new_n479_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1335gat));
  AND4_X1   g505(.A1(new_n240_), .A2(new_n687_), .A3(new_n335_), .A4(new_n683_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n258_), .A3(new_n441_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n651_), .A2(new_n652_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n683_), .A2(new_n240_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n709_), .A2(new_n392_), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n441_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n708_), .B1(new_n713_), .B2(new_n258_), .ZN(G1336gat));
  OAI21_X1  g513(.A(new_n624_), .B1(new_n266_), .B2(new_n265_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT113), .Z(new_n716_));
  NAND2_X1  g515(.A1(new_n711_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n707_), .A2(new_n624_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n260_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT114), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1337gat));
  NAND3_X1  g521(.A1(new_n707_), .A2(new_n283_), .A3(new_n528_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n710_), .A2(new_n392_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n593_), .B(new_n724_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n725_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT115), .B1(new_n725_), .B2(G99gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n707_), .A2(new_n248_), .A3(new_n479_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n479_), .B(new_n724_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(G106gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n731_), .B2(G106gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g535(.A1(new_n392_), .A2(new_n367_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n354_), .A2(new_n356_), .A3(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT12), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n306_), .B2(new_n213_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n351_), .A2(KEYINPUT12), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n321_), .A2(new_n742_), .A3(new_n350_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n743_), .A3(new_n343_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT117), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n345_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n741_), .A2(new_n743_), .A3(KEYINPUT117), .A4(new_n343_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n343_), .A2(new_n345_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT69), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n353_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  AOI22_X1  g550(.A1(new_n746_), .A2(new_n747_), .B1(new_n751_), .B2(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n739_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n365_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(KEYINPUT56), .A3(new_n365_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n737_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n383_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n378_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT118), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT118), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n368_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n659_), .B1(new_n758_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n367_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT56), .B1(new_n753_), .B2(new_n365_), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n755_), .B(new_n364_), .C1(new_n739_), .C2(new_n752_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n772_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n772_), .B(KEYINPUT58), .C1(new_n773_), .C2(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n339_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n737_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n335_), .B1(new_n781_), .B2(new_n766_), .ZN(new_n782_));
  OAI22_X1  g581(.A1(new_n777_), .A2(new_n779_), .B1(new_n782_), .B2(KEYINPUT57), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n770_), .B1(new_n783_), .B2(KEYINPUT120), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n768_), .A2(new_n769_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n775_), .A2(new_n776_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n339_), .A3(new_n778_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n786_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n784_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n240_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n369_), .A2(new_n684_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n341_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n794_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n796_), .A2(new_n241_), .A3(new_n340_), .A4(new_n792_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n791_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n624_), .A2(new_n662_), .A3(new_n529_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n783_), .B2(new_n770_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n782_), .A2(KEYINPUT57), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n785_), .A2(new_n806_), .A3(new_n788_), .A4(KEYINPUT119), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n240_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n799_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(new_n802_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n803_), .B1(new_n810_), .B2(new_n801_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811_), .B2(new_n684_), .ZN(new_n812_));
  INV_X1    g611(.A(G113gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(new_n813_), .A3(new_n392_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1340gat));
  OAI21_X1  g614(.A(G120gat), .B1(new_n811_), .B2(new_n372_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT60), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT121), .B1(new_n817_), .B2(G120gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(G120gat), .B1(new_n683_), .B2(new_n817_), .ZN(new_n819_));
  MUX2_X1   g618(.A(new_n818_), .B(KEYINPUT121), .S(new_n819_), .Z(new_n820_));
  NAND2_X1  g619(.A1(new_n810_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(new_n821_), .ZN(G1341gat));
  OAI21_X1  g621(.A(G127gat), .B1(new_n811_), .B2(new_n240_), .ZN(new_n823_));
  INV_X1    g622(.A(G127gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n810_), .A2(new_n824_), .A3(new_n241_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1342gat));
  OAI21_X1  g625(.A(G134gat), .B1(new_n811_), .B2(new_n340_), .ZN(new_n827_));
  INV_X1    g626(.A(G134gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n810_), .A2(new_n828_), .A3(new_n335_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1343gat));
  NAND3_X1  g629(.A1(new_n785_), .A2(new_n806_), .A3(new_n788_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n241_), .B1(new_n831_), .B2(new_n804_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n798_), .B1(new_n832_), .B2(new_n807_), .ZN(new_n833_));
  OR4_X1    g632(.A1(new_n624_), .A2(new_n833_), .A3(new_n662_), .A4(new_n527_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n684_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT122), .B(G141gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1344gat));
  NOR2_X1   g636(.A1(new_n834_), .A2(new_n372_), .ZN(new_n838_));
  INV_X1    g637(.A(G148gat), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1345gat));
  NOR2_X1   g639(.A1(new_n834_), .A2(new_n240_), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT61), .B(G155gat), .Z(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1346gat));
  OAI21_X1  g642(.A(G162gat), .B1(new_n834_), .B2(new_n340_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n659_), .A2(G162gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n834_), .B2(new_n845_), .ZN(G1347gat));
  AOI21_X1  g645(.A(new_n441_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n848_), .A2(new_n479_), .A3(new_n526_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n241_), .B1(new_n784_), .B2(new_n789_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n392_), .B(new_n849_), .C1(new_n850_), .C2(new_n798_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT62), .B1(new_n851_), .B2(KEYINPUT22), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n800_), .A2(new_n853_), .A3(new_n392_), .A4(new_n849_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n852_), .A2(G169gat), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856_));
  INV_X1    g655(.A(G169gat), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT62), .B(new_n857_), .C1(new_n851_), .C2(KEYINPUT22), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n855_), .A2(new_n856_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n856_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1348gat));
  NOR2_X1   g661(.A1(new_n848_), .A2(new_n526_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(G176gat), .A3(new_n683_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n833_), .A2(new_n864_), .A3(new_n479_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n850_), .A2(new_n798_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n849_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n683_), .ZN(new_n869_));
  INV_X1    g668(.A(G176gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(KEYINPUT124), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(KEYINPUT124), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n865_), .B1(new_n872_), .B2(new_n873_), .ZN(G1349gat));
  NAND2_X1  g673(.A1(new_n241_), .A2(new_n537_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n809_), .A2(new_n241_), .A3(new_n680_), .A4(new_n863_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n868_), .A2(new_n876_), .B1(new_n877_), .B2(new_n487_), .ZN(G1350gat));
  INV_X1    g677(.A(new_n868_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G190gat), .B1(new_n879_), .B2(new_n340_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n868_), .A2(new_n335_), .A3(new_n491_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1351gat));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n847_), .A2(new_n479_), .A3(new_n526_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n833_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n884_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n809_), .A2(KEYINPUT125), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n392_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g689(.A(new_n446_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT125), .B1(new_n809_), .B2(new_n886_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n883_), .B(new_n884_), .C1(new_n808_), .C2(new_n799_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n891_), .B(new_n683_), .C1(new_n892_), .C2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n372_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n894_), .B(new_n895_), .C1(G204gat), .C2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n683_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n899_));
  INV_X1    g698(.A(G204gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n895_), .B1(new_n901_), .B2(new_n894_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n898_), .A2(new_n902_), .ZN(G1353gat));
  NAND2_X1  g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n888_), .A2(new_n241_), .A3(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT127), .ZN(new_n907_));
  XOR2_X1   g706(.A(new_n905_), .B(new_n907_), .Z(G1354gat));
  INV_X1    g707(.A(new_n888_), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n909_), .A2(G218gat), .A3(new_n659_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G218gat), .B1(new_n909_), .B2(new_n340_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1355gat));
endmodule


