//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_;
  XNOR2_X1  g000(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT89), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT90), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n211_), .A3(new_n207_), .A4(new_n208_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n212_), .C1(KEYINPUT1), .C2(new_n203_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT88), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(KEYINPUT88), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n215_), .A2(new_n216_), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT91), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT3), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT91), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n214_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n214_), .B2(new_n220_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT2), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n224_), .A2(new_n226_), .B1(G155gat), .B2(G162gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n207_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n218_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n202_), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n213_), .A2(new_n217_), .B1(new_n227_), .B2(new_n207_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232_));
  INV_X1    g031(.A(new_n202_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G22gat), .B(G50gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n230_), .A2(new_n236_), .A3(new_n234_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT93), .Z(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n232_), .B1(new_n218_), .B2(new_n228_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G211gat), .B(G218gat), .Z(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(G204gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT94), .B(G197gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(G204gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n245_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G204gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n253_), .B(KEYINPUT21), .C1(new_n246_), .C2(new_n252_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n245_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n251_), .A2(new_n254_), .B1(new_n256_), .B2(KEYINPUT21), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n243_), .B1(new_n244_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G78gat), .B(G106gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT95), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n251_), .A2(new_n254_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(KEYINPUT21), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n264_), .B(new_n242_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n261_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n258_), .A2(new_n265_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n259_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n240_), .A2(KEYINPUT96), .A3(new_n266_), .A4(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n268_), .A2(new_n266_), .A3(new_n239_), .A4(new_n238_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT96), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n238_), .A2(new_n239_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n266_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n261_), .B1(new_n258_), .B2(new_n265_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n269_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT27), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT18), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G64gat), .ZN(new_n281_));
  INV_X1    g080(.A(G92gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT98), .A2(G169gat), .A3(G176gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT22), .B(G169gat), .ZN(new_n285_));
  INV_X1    g084(.A(G176gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT98), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n285_), .A2(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(G183gat), .A3(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT84), .ZN(new_n292_));
  INV_X1    g091(.A(G183gat), .ZN(new_n293_));
  INV_X1    g092(.A(G190gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT23), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT84), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(new_n290_), .A3(G183gat), .A4(G190gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n292_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n294_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n298_), .A2(KEYINPUT99), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT99), .B1(new_n298_), .B2(new_n299_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n284_), .B(new_n289_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G169gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n286_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n304_), .A2(KEYINPUT24), .A3(new_n288_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(KEYINPUT24), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n295_), .A2(new_n291_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT26), .B(G190gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT25), .B(G183gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n307_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n302_), .A2(new_n257_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT26), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(G190gat), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n310_), .B(new_n316_), .C1(new_n309_), .C2(new_n314_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n307_), .A2(new_n317_), .A3(new_n298_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n308_), .A2(new_n299_), .ZN(new_n319_));
  OAI21_X1  g118(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n320_));
  OR3_X1    g119(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n264_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n313_), .A2(KEYINPUT20), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT19), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT20), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n302_), .A2(new_n312_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n330_), .B1(new_n331_), .B2(new_n264_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n257_), .A2(new_n322_), .A3(new_n318_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n327_), .B(KEYINPUT97), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n283_), .B1(new_n329_), .B2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n335_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n283_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n339_), .A2(new_n328_), .A3(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n278_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n329_), .A2(new_n337_), .A3(new_n283_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n331_), .A2(new_n264_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n344_), .A2(KEYINPUT20), .A3(new_n333_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n345_), .A2(new_n335_), .B1(new_n327_), .B2(new_n325_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n343_), .B(KEYINPUT27), .C1(new_n346_), .C2(new_n283_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n277_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(KEYINPUT101), .B(KEYINPUT0), .Z(new_n350_));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G57gat), .B(G85gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n356_), .B(KEYINPUT100), .Z(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G127gat), .ZN(new_n359_));
  INV_X1    g158(.A(G134gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G127gat), .A2(G134gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G113gat), .ZN(new_n364_));
  INV_X1    g163(.A(G113gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n365_), .A3(new_n362_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(G120gat), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(G120gat), .B1(new_n364_), .B2(new_n366_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n218_), .A2(new_n370_), .A3(new_n228_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n369_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(KEYINPUT86), .A3(new_n367_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT86), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n218_), .A2(new_n228_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT4), .B1(new_n371_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n373_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n229_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n358_), .B1(new_n377_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n218_), .A2(new_n370_), .A3(new_n228_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n358_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n355_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT4), .B1(new_n229_), .B2(new_n378_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n378_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n383_), .B1(new_n388_), .B2(new_n231_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n389_), .B2(KEYINPUT4), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n354_), .B(new_n384_), .C1(new_n390_), .C2(new_n358_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT85), .B(KEYINPUT30), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n378_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G71gat), .B(G99gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G15gat), .B(G43gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT31), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(new_n323_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n397_), .B(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n349_), .A2(new_n393_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT105), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT105), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n349_), .A2(new_n406_), .A3(new_n393_), .A4(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n283_), .A2(KEYINPUT32), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n346_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n329_), .A2(new_n337_), .A3(new_n409_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT103), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT103), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n329_), .A2(new_n337_), .A3(new_n413_), .A4(new_n409_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n392_), .A2(new_n410_), .A3(new_n412_), .A4(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n338_), .A2(new_n341_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n391_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n377_), .A2(new_n381_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n357_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n420_), .A2(KEYINPUT33), .A3(new_n354_), .A4(new_n384_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT102), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n389_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n379_), .A2(KEYINPUT102), .A3(new_n383_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n357_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n425_), .B(new_n355_), .C1(new_n357_), .C2(new_n390_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n416_), .A2(new_n418_), .A3(new_n421_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n415_), .A2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n269_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n428_), .A2(KEYINPUT104), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT104), .B1(new_n428_), .B2(new_n429_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n429_), .A2(new_n392_), .A3(new_n348_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n403_), .B(KEYINPUT87), .Z(new_n434_));
  OAI21_X1  g233(.A(new_n408_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(G230gat), .A2(G233gat), .ZN(new_n436_));
  INV_X1    g235(.A(G99gat), .ZN(new_n437_));
  INV_X1    g236(.A(G106gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT65), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n437_), .B(new_n438_), .C1(new_n439_), .C2(KEYINPUT7), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT7), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n441_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT67), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT66), .ZN(new_n446_));
  NAND3_X1  g245(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n446_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G99gat), .A2(G106gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(KEYINPUT66), .A3(new_n447_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT67), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n445_), .A2(new_n450_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G85gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n282_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT8), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n460_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(KEYINPUT8), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n458_), .A2(KEYINPUT9), .A3(new_n459_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n459_), .A2(KEYINPUT9), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT10), .B(G99gat), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n467_), .B(new_n468_), .C1(G106gat), .C2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n443_), .A2(new_n461_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n453_), .A2(KEYINPUT64), .A3(new_n447_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n472_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n463_), .A2(new_n466_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT68), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT68), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n463_), .A2(new_n478_), .A3(new_n481_), .A4(new_n466_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n485_));
  XOR2_X1   g284(.A(G71gat), .B(G78gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n436_), .B1(new_n483_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n479_), .A2(KEYINPUT12), .A3(new_n489_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n480_), .A2(new_n482_), .A3(new_n489_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n494_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n491_), .B(new_n492_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT69), .B1(new_n483_), .B2(new_n490_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n501_));
  AOI211_X1 g300(.A(new_n501_), .B(new_n489_), .C1(new_n480_), .C2(new_n482_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT70), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n462_), .A2(new_n456_), .B1(new_n472_), .B2(new_n477_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n481_), .B1(new_n504_), .B2(new_n466_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n462_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT67), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT67), .B1(new_n440_), .B2(new_n442_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n450_), .A2(new_n454_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n506_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n476_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n512_));
  NOR4_X1   g311(.A1(new_n511_), .A2(new_n512_), .A3(KEYINPUT68), .A4(new_n465_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n490_), .B1(new_n505_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n501_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT70), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n483_), .A2(KEYINPUT69), .A3(new_n490_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n503_), .A2(new_n518_), .A3(new_n493_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n499_), .B1(new_n436_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G120gat), .B(G148gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT5), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G176gat), .B(G204gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  NOR2_X1   g325(.A1(new_n520_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n519_), .A2(new_n436_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n498_), .A3(new_n526_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(KEYINPUT13), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT13), .ZN(new_n532_));
  INV_X1    g331(.A(new_n530_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n532_), .B1(new_n527_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(new_n303_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n246_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(G50gat), .ZN(new_n540_));
  OR2_X1    g339(.A1(G29gat), .A2(G36gat), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT76), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n542_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n545_), .A2(G43gat), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(G43gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G29gat), .B(G36gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT76), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n550_), .B2(new_n544_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n540_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(G43gat), .B1(new_n545_), .B2(new_n546_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n550_), .A2(new_n548_), .A3(new_n544_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(G50gat), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G1gat), .ZN(new_n557_));
  INV_X1    g356(.A(G8gat), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT14), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT79), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT79), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n562_), .B(KEYINPUT14), .C1(new_n557_), .C2(new_n558_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G1gat), .B(G8gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n556_), .A2(KEYINPUT81), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT81), .B1(new_n556_), .B2(new_n566_), .ZN(new_n569_));
  OAI22_X1  g368(.A1(new_n568_), .A2(new_n569_), .B1(new_n566_), .B2(new_n556_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(G229gat), .A3(G233gat), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT15), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n547_), .A2(new_n551_), .A3(new_n540_), .ZN(new_n573_));
  AOI21_X1  g372(.A(G50gat), .B1(new_n553_), .B2(new_n554_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n566_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n552_), .A2(KEYINPUT15), .A3(new_n555_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT82), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n578_), .B(new_n581_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n539_), .B1(new_n571_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n556_), .A2(new_n566_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT81), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n556_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n586_), .A2(new_n567_), .B1(new_n576_), .B2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n582_), .B(new_n539_), .C1(new_n588_), .C2(new_n579_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n583_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n535_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n435_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT16), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(G183gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G211gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n489_), .B(new_n566_), .Z(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n597_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT17), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n601_), .A2(new_n597_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT77), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n556_), .B1(new_n505_), .B2(new_n513_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n575_), .A2(new_n577_), .A3(new_n479_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT75), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n608_), .B1(new_n611_), .B2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n587_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n575_), .A2(new_n577_), .A3(new_n479_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n608_), .B(new_n616_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT36), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n360_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(G162gat), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n618_), .A2(new_n619_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n614_), .A2(new_n615_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n616_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n622_), .A2(new_n623_), .A3(new_n626_), .A4(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT78), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT77), .B1(new_n627_), .B2(new_n629_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n630_), .A3(new_n620_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n626_), .A2(new_n623_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n626_), .A2(new_n623_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n631_), .A2(new_n632_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT37), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n631_), .A2(new_n637_), .A3(new_n632_), .A4(KEYINPUT37), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n593_), .A2(new_n607_), .A3(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n557_), .A3(new_n392_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT38), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n631_), .A2(new_n637_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT106), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n593_), .A2(new_n647_), .A3(new_n607_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(new_n392_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n557_), .B2(new_n649_), .ZN(G1324gat));
  AOI21_X1  g449(.A(new_n558_), .B1(new_n648_), .B2(new_n348_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT39), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n643_), .A2(new_n558_), .A3(new_n348_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1325gat));
  INV_X1    g455(.A(G15gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n648_), .B2(new_n434_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT41), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n643_), .A2(new_n657_), .A3(new_n434_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1326gat));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n648_), .B2(new_n277_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT42), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n643_), .A2(new_n662_), .A3(new_n277_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n435_), .A2(new_n642_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT43), .B1(new_n667_), .B2(KEYINPUT107), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n669_), .B(new_n670_), .C1(new_n435_), .C2(new_n642_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n592_), .B(new_n607_), .C1(new_n668_), .C2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n428_), .A2(new_n429_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n429_), .A2(new_n348_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n393_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n428_), .A2(KEYINPUT104), .A3(new_n429_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n434_), .ZN(new_n682_));
  AOI22_X1  g481(.A1(new_n681_), .A2(new_n682_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n640_), .A2(new_n641_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n670_), .B1(new_n685_), .B2(new_n669_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n667_), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n688_), .A2(KEYINPUT44), .A3(new_n592_), .A4(new_n607_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n674_), .A2(new_n392_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G29gat), .ZN(new_n691_));
  INV_X1    g490(.A(new_n646_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n593_), .A2(new_n692_), .A3(new_n606_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n393_), .A2(G29gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n606_), .A2(new_n692_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n435_), .A2(new_n592_), .A3(new_n698_), .A4(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n348_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT108), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n700_), .A2(KEYINPUT108), .A3(new_n701_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n697_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n704_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(KEYINPUT45), .A3(new_n702_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n674_), .A2(new_n348_), .A3(new_n689_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(G36gat), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n712_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n710_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n713_), .A2(new_n716_), .ZN(G1329gat));
  NAND3_X1  g516(.A1(new_n674_), .A2(new_n403_), .A3(new_n689_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G43gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n693_), .A2(new_n548_), .A3(new_n434_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(G1330gat));
  NAND3_X1  g522(.A1(new_n674_), .A2(new_n277_), .A3(new_n689_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n725_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(G50gat), .A3(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n693_), .A2(new_n540_), .A3(new_n277_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1331gat));
  INV_X1    g529(.A(new_n591_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n535_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n683_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n607_), .A2(new_n642_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n392_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n732_), .A2(new_n731_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n435_), .A2(new_n737_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n738_), .A2(new_n647_), .A3(new_n607_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n392_), .A2(G57gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1332gat));
  INV_X1    g540(.A(G64gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n739_), .B2(new_n348_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT48), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n735_), .A2(new_n742_), .A3(new_n348_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n739_), .B2(new_n434_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT49), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n735_), .A2(new_n747_), .A3(new_n434_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n739_), .B2(new_n277_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT50), .Z(new_n754_));
  NAND3_X1  g553(.A1(new_n735_), .A2(new_n752_), .A3(new_n277_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n738_), .A2(new_n692_), .A3(new_n606_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n392_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n737_), .A2(new_n607_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n393_), .A2(new_n457_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n758_), .B1(new_n760_), .B2(new_n761_), .ZN(G1336gat));
  AOI21_X1  g561(.A(G92gat), .B1(new_n757_), .B2(new_n348_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n701_), .A2(new_n282_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n760_), .B2(new_n764_), .ZN(G1337gat));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n437_), .B1(new_n760_), .B2(new_n434_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769_));
  INV_X1    g568(.A(new_n469_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n757_), .A2(new_n770_), .A3(new_n403_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n769_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n769_), .B1(new_n768_), .B2(new_n771_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n766_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n774_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(KEYINPUT51), .A3(new_n772_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1338gat));
  AOI211_X1 g577(.A(new_n429_), .B(new_n759_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT114), .B1(new_n779_), .B2(new_n438_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n760_), .A2(new_n277_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(G106gat), .ZN(new_n783_));
  XOR2_X1   g582(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n757_), .A2(new_n438_), .A3(new_n277_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT112), .Z(new_n787_));
  INV_X1    g586(.A(new_n784_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT114), .B(new_n788_), .C1(new_n779_), .C2(new_n438_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT53), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n785_), .A2(new_n787_), .A3(new_n792_), .A4(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1339gat));
  NAND4_X1  g593(.A1(new_n732_), .A2(KEYINPUT54), .A3(new_n591_), .A4(new_n734_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n684_), .A2(new_n591_), .A3(new_n606_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n535_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n795_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n492_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n500_), .A2(new_n502_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n436_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n498_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n493_), .A2(new_n495_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT72), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n808_), .A2(KEYINPUT55), .A3(new_n491_), .A4(new_n492_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n802_), .A2(new_n804_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n526_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(new_n814_), .A3(new_n811_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n578_), .B(new_n580_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n538_), .C1(new_n588_), .C2(new_n580_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n589_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT116), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n589_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n530_), .A2(KEYINPUT118), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT118), .B1(new_n530_), .B2(new_n822_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n813_), .B(new_n815_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT119), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n684_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n814_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n530_), .A2(new_n822_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n530_), .A2(KEYINPUT118), .A3(new_n822_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n829_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(KEYINPUT58), .A4(new_n815_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n827_), .A2(new_n828_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n822_), .B1(new_n527_), .B2(new_n533_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n591_), .B1(new_n520_), .B2(new_n526_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n841_), .B2(KEYINPUT56), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n840_), .B(new_n814_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n692_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n844_), .A2(new_n692_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n845_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n837_), .A2(new_n847_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n799_), .B1(new_n850_), .B2(new_n607_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n349_), .A2(new_n392_), .A3(new_n403_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT120), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT59), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n812_), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n839_), .C1(KEYINPUT56), .C2(new_n841_), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n646_), .B(new_n845_), .C1(new_n858_), .C2(new_n838_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n846_), .B1(new_n844_), .B2(new_n692_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n606_), .B1(new_n861_), .B2(new_n837_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n856_), .B(new_n853_), .C1(new_n862_), .C2(new_n799_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n855_), .A2(new_n731_), .A3(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n851_), .A2(new_n854_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n591_), .A2(G113gat), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n864_), .A2(G113gat), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT121), .ZN(G1340gat));
  NAND3_X1  g667(.A1(new_n855_), .A2(new_n535_), .A3(new_n863_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n855_), .A2(new_n863_), .A3(KEYINPUT122), .A4(new_n535_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(G120gat), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n732_), .B2(G120gat), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n865_), .B(new_n875_), .C1(new_n874_), .C2(G120gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT123), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n873_), .A2(new_n879_), .A3(new_n876_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1341gat));
  AOI21_X1  g680(.A(G127gat), .B1(new_n865_), .B2(new_n606_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n855_), .A2(new_n863_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n607_), .A2(new_n359_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1342gat));
  AOI21_X1  g684(.A(G134gat), .B1(new_n865_), .B2(new_n647_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n684_), .A2(new_n360_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n883_), .B2(new_n887_), .ZN(G1343gat));
  NOR2_X1   g687(.A1(new_n851_), .A2(new_n434_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n392_), .A3(new_n678_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT124), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n889_), .A2(new_n892_), .A3(new_n392_), .A4(new_n678_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n591_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(G141gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1344gat));
  AOI21_X1  g695(.A(new_n732_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n897_));
  INV_X1    g696(.A(G148gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1345gat));
  AOI21_X1  g698(.A(new_n607_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT61), .B(G155gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  NAND2_X1  g701(.A1(new_n891_), .A2(new_n893_), .ZN(new_n903_));
  AOI21_X1  g702(.A(G162gat), .B1(new_n903_), .B2(new_n647_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n684_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(G162gat), .B2(new_n905_), .ZN(G1347gat));
  NOR3_X1   g705(.A1(new_n701_), .A2(new_n277_), .A3(new_n392_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n434_), .B(new_n907_), .C1(new_n862_), .C2(new_n799_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n591_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n909_), .A2(new_n285_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n303_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT62), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(KEYINPUT62), .B2(new_n911_), .ZN(G1348gat));
  NOR2_X1   g712(.A1(new_n908_), .A2(new_n732_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n286_), .ZN(G1349gat));
  NOR2_X1   g714(.A1(new_n908_), .A2(new_n607_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n310_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n293_), .B2(new_n916_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n908_), .B2(new_n684_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n647_), .A2(new_n309_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n908_), .B2(new_n920_), .ZN(G1351gat));
  NOR3_X1   g720(.A1(new_n429_), .A2(new_n701_), .A3(new_n392_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n889_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n591_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n246_), .ZN(G1352gat));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n732_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n252_), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT125), .B(G204gat), .Z(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n926_), .B2(new_n929_), .ZN(G1353gat));
  NOR2_X1   g729(.A1(new_n923_), .A2(new_n607_), .ZN(new_n931_));
  OR2_X1    g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n931_), .A2(new_n932_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(G1354gat));
  INV_X1    g737(.A(new_n923_), .ZN(new_n939_));
  AOI21_X1  g738(.A(G218gat), .B1(new_n939_), .B2(new_n647_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n642_), .A2(G218gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT127), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n939_), .B2(new_n942_), .ZN(G1355gat));
endmodule


