//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT64), .B1(G85gat), .B2(G92gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n214_), .B(new_n217_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n216_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n225_), .A2(new_n212_), .A3(new_n213_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  XOR2_X1   g027(.A(G85gat), .B(G92gat), .Z(new_n229_));
  AND3_X1   g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n222_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n209_), .A2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n208_), .B(new_n222_), .C1(new_n231_), .C2(new_n230_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(KEYINPUT12), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT12), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n209_), .A2(new_n232_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G230gat), .A2(G233gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n233_), .A2(new_n234_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n239_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G120gat), .B(G148gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G204gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT5), .B(G176gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n240_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n248_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT13), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n254_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G113gat), .B(G141gat), .ZN(new_n259_));
  INV_X1    g058(.A(G197gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT72), .B(G169gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G1gat), .ZN(new_n265_));
  INV_X1    g064(.A(G8gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT14), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G15gat), .B(G22gat), .ZN(new_n270_));
  OAI211_X1 g069(.A(KEYINPUT68), .B(KEYINPUT14), .C1(new_n265_), .C2(new_n266_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G1gat), .B(G8gat), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n269_), .A2(new_n273_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT66), .B(G29gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G43gat), .B(G50gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(G36gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n280_), .A2(G36gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n279_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n280_), .A2(G36gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(new_n278_), .A3(new_n281_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n284_), .A2(KEYINPUT15), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT15), .B1(new_n284_), .B2(new_n286_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n277_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G229gat), .A2(G233gat), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n284_), .A2(new_n286_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n284_), .A2(new_n286_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(KEYINPUT71), .A3(new_n291_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n297_));
  INV_X1    g096(.A(new_n291_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n297_), .B1(new_n298_), .B2(new_n294_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n290_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n264_), .B1(new_n293_), .B2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n290_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n304_), .A2(new_n292_), .A3(new_n263_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n258_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G190gat), .B(G218gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G134gat), .B(G162gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(KEYINPUT36), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n284_), .A2(new_n286_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n232_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT67), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G232gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT34), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n318_), .A2(KEYINPUT35), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n232_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n316_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(KEYINPUT35), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n316_), .A2(new_n320_), .A3(KEYINPUT35), .A4(new_n318_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n313_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n322_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n313_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n311_), .A2(new_n312_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n327_), .B(new_n324_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G183gat), .A3(G190gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(G190gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT23), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n332_), .A2(KEYINPUT76), .A3(G183gat), .A4(G190gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(KEYINPUT75), .A2(G169gat), .A3(G176gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n341_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT77), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT25), .B(G183gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT26), .B1(new_n349_), .B2(new_n337_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT26), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT74), .A3(G190gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n348_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354_));
  INV_X1    g153(.A(G169gat), .ZN(new_n355_));
  INV_X1    g154(.A(G176gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n357_), .A2(KEYINPUT24), .A3(new_n358_), .A4(new_n342_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n340_), .A2(new_n361_), .A3(new_n345_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n347_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n338_), .A2(new_n333_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n336_), .A2(new_n337_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n355_), .B2(KEYINPUT22), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT22), .B(G169gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n367_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT79), .B(G176gat), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n366_), .B(new_n358_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n363_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n260_), .A3(G204gat), .ZN(new_n375_));
  INV_X1    g174(.A(G204gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT87), .B1(new_n376_), .B2(G197gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(G197gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n375_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G211gat), .B(G218gat), .Z(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(KEYINPUT21), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT88), .ZN(new_n382_));
  INV_X1    g181(.A(new_n380_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n260_), .A2(G204gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT21), .B1(new_n378_), .B2(new_n384_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n383_), .B(new_n385_), .C1(new_n379_), .C2(KEYINPUT21), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n379_), .A2(new_n387_), .A3(KEYINPUT21), .A4(new_n380_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n373_), .A2(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n382_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n371_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n369_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n358_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n340_), .A2(KEYINPUT92), .A3(new_n365_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT92), .B1(new_n340_), .B2(new_n365_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n395_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n400_));
  AND2_X1   g199(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n401_));
  AND2_X1   g200(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n403_));
  OAI22_X1  g202(.A1(new_n400_), .A2(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n345_), .A2(new_n359_), .A3(new_n364_), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT91), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT26), .B(G190gat), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n348_), .A2(new_n407_), .B1(new_n338_), .B2(new_n333_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n359_), .A4(new_n345_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n391_), .A2(new_n399_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n413_), .B(KEYINPUT19), .Z(new_n414_));
  NAND4_X1  g213(.A1(new_n390_), .A2(KEYINPUT20), .A3(new_n412_), .A4(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT93), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n406_), .A2(new_n410_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n340_), .A2(new_n365_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT92), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n394_), .B1(new_n420_), .B2(new_n396_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n389_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n391_), .A2(new_n372_), .A3(new_n363_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(KEYINPUT20), .A3(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n414_), .B(KEYINPUT90), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n373_), .B2(new_n389_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT93), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n414_), .A4(new_n412_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n416_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G92gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT18), .B(G64gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n416_), .A2(new_n427_), .A3(new_n436_), .A4(new_n431_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT27), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n422_), .A2(KEYINPUT20), .A3(new_n425_), .A4(new_n423_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT97), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n399_), .A2(new_n411_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n428_), .B1(new_n444_), .B2(new_n389_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT97), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n425_), .A4(new_n423_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n399_), .A2(new_n405_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT96), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT96), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n399_), .A2(new_n451_), .A3(new_n405_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n391_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n414_), .B1(new_n453_), .B2(new_n429_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n436_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n439_), .A2(KEYINPUT27), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n456_), .A2(KEYINPUT99), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT99), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n439_), .A2(KEYINPUT27), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n443_), .A2(new_n447_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n437_), .B1(new_n461_), .B2(new_n454_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n459_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n441_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT100), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G127gat), .B(G134gat), .ZN(new_n467_));
  INV_X1    g266(.A(G120gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT82), .B(G113gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT30), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n373_), .B(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT81), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT31), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G71gat), .B(G99gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT80), .ZN(new_n479_));
  XOR2_X1   g278(.A(G15gat), .B(G43gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G227gat), .A2(G233gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  NAND3_X1  g282(.A1(new_n476_), .A2(new_n477_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n477_), .B1(new_n476_), .B2(new_n483_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n472_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n476_), .A2(new_n483_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT31), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(new_n471_), .A3(new_n484_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n474_), .A2(new_n475_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n487_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(G155gat), .A2(G162gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n494_), .B(KEYINPUT83), .Z(new_n495_));
  NAND2_X1  g294(.A1(G155gat), .A2(G162gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT3), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT2), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G141gat), .A2(G148gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n499_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n500_), .B2(new_n499_), .ZN(new_n503_));
  OAI221_X1 g302(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n497_), .A2(KEYINPUT3), .ZN(new_n505_));
  INV_X1    g304(.A(G141gat), .ZN(new_n506_));
  INV_X1    g305(.A(G148gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n505_), .B(new_n508_), .Z(new_n509_));
  OAI211_X1 g308(.A(new_n495_), .B(new_n496_), .C1(new_n504_), .C2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n496_), .B(KEYINPUT1), .Z(new_n511_));
  NAND2_X1  g310(.A1(new_n495_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n508_), .A3(new_n500_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n472_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n471_), .A2(new_n513_), .A3(new_n510_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(KEYINPUT4), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G225gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT4), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n472_), .A2(new_n520_), .A3(new_n514_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n515_), .A2(new_n518_), .A3(new_n516_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G29gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT95), .ZN(new_n526_));
  XOR2_X1   g325(.A(G57gat), .B(G85gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n524_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n522_), .A2(new_n523_), .A3(new_n530_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n492_), .A2(new_n493_), .A3(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT100), .B(new_n441_), .C1(new_n458_), .C2(new_n463_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n391_), .B1(new_n514_), .B2(KEYINPUT29), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G228gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G78gat), .B(G106gat), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n514_), .A2(KEYINPUT29), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n544_));
  XNOR2_X1  g343(.A(G22gat), .B(G50gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n543_), .B(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT89), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n539_), .A2(new_n541_), .ZN(new_n549_));
  OR3_X1    g348(.A1(new_n542_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n547_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n542_), .A2(KEYINPUT89), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n466_), .A2(new_n535_), .A3(new_n536_), .A4(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n493_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n487_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n533_), .B(KEYINPUT33), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n517_), .A2(new_n518_), .A3(new_n521_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n515_), .A2(new_n519_), .A3(new_n516_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n531_), .A3(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n558_), .A2(new_n439_), .A3(new_n438_), .A4(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n436_), .A2(KEYINPUT32), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n461_), .B2(new_n454_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT98), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n432_), .A2(new_n563_), .ZN(new_n567_));
  OAI211_X1 g366(.A(KEYINPUT98), .B(new_n563_), .C1(new_n461_), .C2(new_n454_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n566_), .A2(new_n534_), .A3(new_n567_), .A4(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n562_), .A2(new_n553_), .A3(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT99), .B1(new_n456_), .B2(new_n457_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n460_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n534_), .B(new_n440_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n557_), .B(new_n570_), .C1(new_n573_), .C2(new_n553_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n331_), .B1(new_n554_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n208_), .B(new_n277_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT69), .B(KEYINPUT16), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G127gat), .B(G155gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n583_), .A2(new_n584_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n578_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n585_), .B2(new_n578_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT70), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n308_), .A2(new_n575_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n534_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n258_), .B1(new_n554_), .B2(new_n574_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n331_), .A2(KEYINPUT37), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n326_), .A2(new_n596_), .A3(new_n330_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(new_n589_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n306_), .B(KEYINPUT73), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n594_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n534_), .B(KEYINPUT101), .Z(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n265_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT102), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n605_), .A2(KEYINPUT38), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(KEYINPUT38), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n593_), .B1(new_n606_), .B2(new_n607_), .ZN(G1324gat));
  NAND2_X1  g407(.A1(new_n466_), .A2(new_n536_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n602_), .A2(new_n266_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G8gat), .B1(new_n591_), .B2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(KEYINPUT39), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(KEYINPUT39), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n610_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g415(.A(G15gat), .B1(new_n591_), .B2(new_n557_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT41), .Z(new_n618_));
  INV_X1    g417(.A(G15gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n557_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n602_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n621_), .ZN(G1326gat));
  NOR2_X1   g421(.A1(new_n553_), .A2(G22gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT104), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n602_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G22gat), .B1(new_n591_), .B2(new_n553_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT103), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT42), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n629_), .B(G22gat), .C1(new_n591_), .C2(new_n553_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n627_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n625_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(KEYINPUT105), .B(new_n625_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1327gat));
  NAND2_X1  g436(.A1(new_n589_), .A2(new_n331_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT107), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n594_), .A2(new_n601_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(G29gat), .B1(new_n640_), .B2(new_n534_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n598_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n554_), .A2(new_n574_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(new_n598_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n598_), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n648_), .B(new_n644_), .C1(new_n554_), .C2(new_n574_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n589_), .B(new_n308_), .C1(new_n647_), .C2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n652_), .A2(G29gat), .A3(new_n603_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n648_), .B1(new_n554_), .B2(new_n574_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(new_n645_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n655_), .A2(KEYINPUT44), .A3(new_n589_), .A4(new_n308_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n641_), .B1(new_n653_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658_));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n640_), .A2(KEYINPUT45), .A3(new_n659_), .A4(new_n609_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT45), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n594_), .A2(new_n659_), .A3(new_n601_), .A4(new_n639_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(new_n611_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n656_), .A2(new_n652_), .A3(new_n609_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(G36gat), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n658_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n611_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n659_), .B1(new_n669_), .B2(new_n656_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT108), .B(KEYINPUT46), .C1(new_n670_), .C2(new_n664_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n668_), .A2(new_n671_), .ZN(G1329gat));
  NAND4_X1  g471(.A1(new_n656_), .A2(new_n652_), .A3(G43gat), .A4(new_n620_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n640_), .A2(new_n620_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(G43gat), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g475(.A(new_n553_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G50gat), .B1(new_n640_), .B2(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n656_), .A2(new_n652_), .A3(G50gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(new_n677_), .ZN(G1331gat));
  NOR2_X1   g479(.A1(new_n257_), .A2(new_n589_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n575_), .A2(new_n600_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n592_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n258_), .A2(new_n599_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT109), .Z(new_n686_));
  AOI21_X1  g485(.A(new_n306_), .B1(new_n554_), .B2(new_n574_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n603_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n684_), .B1(new_n689_), .B2(new_n683_), .ZN(G1332gat));
  INV_X1    g489(.A(G64gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n691_), .A3(new_n609_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G64gat), .B1(new_n682_), .B2(new_n611_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(KEYINPUT48), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n693_), .A2(KEYINPUT48), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n692_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT110), .ZN(G1333gat));
  INV_X1    g496(.A(G71gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n688_), .A2(new_n698_), .A3(new_n620_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n682_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n700_), .B2(new_n620_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT49), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n702_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n699_), .B1(new_n706_), .B2(new_n707_), .ZN(G1334gat));
  INV_X1    g507(.A(G78gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n688_), .A2(new_n709_), .A3(new_n677_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G78gat), .B1(new_n682_), .B2(new_n553_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT50), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1335gat));
  AND3_X1   g512(.A1(new_n687_), .A2(new_n258_), .A3(new_n639_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n603_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n257_), .A2(new_n590_), .A3(new_n306_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n655_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n534_), .A2(G85gat), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT112), .Z(new_n719_));
  AOI21_X1  g518(.A(new_n715_), .B1(new_n717_), .B2(new_n719_), .ZN(G1336gat));
  AOI21_X1  g519(.A(G92gat), .B1(new_n714_), .B2(new_n609_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n609_), .A2(G92gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n717_), .B2(new_n722_), .ZN(G1337gat));
  AOI21_X1  g522(.A(new_n224_), .B1(new_n717_), .B2(new_n620_), .ZN(new_n724_));
  AND2_X1   g523(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n714_), .A2(new_n620_), .A3(new_n215_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(G1338gat));
  NAND4_X1  g528(.A1(new_n655_), .A2(KEYINPUT115), .A3(new_n677_), .A4(new_n716_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n677_), .B(new_n716_), .C1(new_n647_), .C2(new_n649_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n733_), .A3(G106gat), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n730_), .A2(new_n733_), .A3(KEYINPUT52), .A4(G106gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n714_), .A2(new_n216_), .A3(new_n677_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT114), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n737_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT53), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n736_), .A2(new_n742_), .A3(new_n737_), .A4(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1339gat));
  INV_X1    g543(.A(new_n253_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n599_), .A2(new_n745_), .A3(new_n600_), .A4(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n240_), .A2(KEYINPUT118), .A3(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n235_), .A2(new_n242_), .A3(new_n237_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n242_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT118), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT55), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n751_), .A2(new_n752_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n247_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT119), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n247_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n249_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT117), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n756_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n247_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n763_), .A2(KEYINPUT117), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n762_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n289_), .A2(new_n301_), .A3(new_n291_), .ZN(new_n769_));
  AOI211_X1 g568(.A(new_n264_), .B(new_n769_), .C1(new_n290_), .C2(new_n300_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n770_), .A2(new_n305_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(new_n252_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n331_), .B1(new_n768_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT122), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT57), .B1(new_n773_), .B2(KEYINPUT122), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n771_), .A2(new_n250_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n759_), .B(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n761_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT58), .B(new_n778_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n598_), .A3(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT122), .B(KEYINPUT57), .C1(new_n773_), .C2(new_n774_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n777_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n749_), .B1(new_n788_), .B2(new_n589_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n609_), .A2(new_n677_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n790_), .A2(new_n603_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT123), .B1(new_n791_), .B2(new_n620_), .ZN(new_n792_));
  AND4_X1   g591(.A1(KEYINPUT123), .A2(new_n790_), .A3(new_n620_), .A4(new_n603_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n789_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G113gat), .B1(new_n794_), .B2(new_n306_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n789_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT125), .B1(new_n792_), .B2(new_n793_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(KEYINPUT124), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT124), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT125), .B1(new_n801_), .B2(new_n799_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n794_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n600_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n795_), .B1(new_n804_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g604(.A(new_n468_), .B1(new_n257_), .B2(KEYINPUT60), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n794_), .B(new_n806_), .C1(KEYINPUT60), .C2(new_n468_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n257_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n468_), .ZN(G1341gat));
  AOI21_X1  g608(.A(G127gat), .B1(new_n794_), .B2(new_n590_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n589_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g611(.A(G134gat), .B1(new_n794_), .B2(new_n331_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n648_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(G134gat), .ZN(G1343gat));
  NOR4_X1   g614(.A1(new_n789_), .A2(new_n609_), .A3(new_n553_), .A4(new_n620_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n603_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n506_), .A3(new_n306_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G141gat), .B1(new_n817_), .B2(new_n307_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1344gat));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n507_), .A3(new_n258_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G148gat), .B1(new_n817_), .B2(new_n257_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1345gat));
  XNOR2_X1  g623(.A(KEYINPUT61), .B(G155gat), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n817_), .B2(new_n589_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n816_), .A2(new_n590_), .A3(new_n603_), .A4(new_n825_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1346gat));
  INV_X1    g628(.A(G162gat), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n648_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n816_), .A2(new_n331_), .A3(new_n603_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n818_), .A2(new_n831_), .B1(new_n832_), .B2(new_n830_), .ZN(G1347gat));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n611_), .A2(new_n603_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n557_), .A2(new_n677_), .ZN(new_n836_));
  AND4_X1   g635(.A1(new_n306_), .A2(new_n796_), .A3(new_n835_), .A4(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n834_), .B1(new_n837_), .B2(new_n355_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n789_), .A2(new_n677_), .A3(new_n557_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n835_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT62), .B(G169gat), .C1(new_n840_), .C2(new_n307_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n369_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(new_n841_), .A3(new_n842_), .ZN(G1348gat));
  NOR3_X1   g642(.A1(new_n840_), .A2(new_n356_), .A3(new_n257_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n840_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n258_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n392_), .B2(new_n846_), .ZN(G1349gat));
  NOR2_X1   g646(.A1(new_n840_), .A2(new_n589_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n348_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n336_), .B2(new_n848_), .ZN(G1350gat));
  OAI21_X1  g649(.A(G190gat), .B1(new_n840_), .B2(new_n648_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n331_), .A2(new_n407_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n840_), .B2(new_n852_), .ZN(G1351gat));
  NOR3_X1   g652(.A1(new_n789_), .A2(new_n553_), .A3(new_n620_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n611_), .A2(new_n534_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(new_n260_), .A3(new_n306_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G197gat), .B1(new_n856_), .B2(new_n307_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1352gat));
  NOR2_X1   g659(.A1(new_n856_), .A2(new_n257_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT126), .B(G204gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n861_), .B2(new_n864_), .ZN(G1353gat));
  NAND3_X1  g664(.A1(new_n854_), .A2(new_n590_), .A3(new_n855_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT63), .B(G211gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n866_), .B2(new_n869_), .ZN(G1354gat));
  NAND2_X1  g669(.A1(new_n788_), .A2(new_n589_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n749_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n553_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n873_), .A2(new_n557_), .A3(new_n331_), .A4(new_n855_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT127), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n854_), .A2(KEYINPUT127), .A3(new_n331_), .A4(new_n855_), .ZN(new_n877_));
  INV_X1    g676(.A(G218gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n857_), .A2(G218gat), .A3(new_n598_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1355gat));
endmodule


