//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  AND3_X1   g007(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n203_), .A2(new_n204_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n208_), .A2(new_n211_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT95), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT22), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G169gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n206_), .A2(KEYINPUT22), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n207_), .ZN(new_n221_));
  AND3_X1   g020(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT94), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n222_), .A2(new_n223_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT94), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n220_), .A3(new_n207_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n209_), .A2(new_n210_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n217_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n234_));
  AOI211_X1 g033(.A(KEYINPUT95), .B(new_n232_), .C1(new_n225_), .C2(new_n229_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n216_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT87), .B(G197gat), .ZN(new_n238_));
  OAI211_X1 g037(.A(KEYINPUT21), .B(new_n237_), .C1(new_n238_), .C2(G204gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(G211gat), .B(G218gat), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G197gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT88), .B1(new_n242_), .B2(G204gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT88), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(G197gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n245_), .B2(new_n238_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n239_), .B(new_n241_), .C1(new_n248_), .C2(KEYINPUT21), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n242_), .A2(KEYINPUT87), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT87), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G197gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n253_), .A2(G204gat), .B1(new_n243_), .B2(new_n246_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n240_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n247_), .B(new_n255_), .C1(new_n245_), .C2(new_n238_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT21), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n249_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n236_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G183gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT75), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT75), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(G183gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n264_), .A3(KEYINPUT25), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT76), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n261_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT75), .B(G183gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT76), .B1(new_n270_), .B2(new_n267_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n271_), .A3(new_n212_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n204_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n273_), .A2(KEYINPUT24), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n272_), .A2(new_n274_), .A3(new_n211_), .A4(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n211_), .B1(G190gat), .B2(new_n270_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT78), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n220_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n206_), .A2(KEYINPUT78), .A3(KEYINPUT22), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n207_), .A4(new_n219_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n226_), .A3(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT90), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n259_), .A2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n243_), .A2(new_n246_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n245_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT89), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n288_), .A2(KEYINPUT21), .A3(new_n240_), .A4(new_n257_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(KEYINPUT90), .A3(new_n249_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n283_), .A2(new_n285_), .A3(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n260_), .A2(new_n291_), .A3(KEYINPUT20), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT19), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296_));
  INV_X1    g095(.A(G92gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT18), .B(G64gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n259_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n302_), .B(new_n216_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n276_), .A2(new_n282_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n289_), .A2(KEYINPUT90), .A3(new_n249_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT90), .B1(new_n289_), .B2(new_n249_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n294_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n303_), .A2(new_n307_), .A3(KEYINPUT20), .A4(new_n308_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n295_), .A2(new_n301_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n230_), .A2(new_n233_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n302_), .A2(new_n216_), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n307_), .A2(KEYINPUT20), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n294_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n260_), .A2(new_n291_), .A3(KEYINPUT20), .A4(new_n308_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n301_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n310_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT20), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n305_), .A2(new_n306_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n320_), .B2(new_n283_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n308_), .B1(new_n321_), .B2(new_n260_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n309_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n300_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n295_), .A2(new_n301_), .A3(new_n309_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT27), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n202_), .B1(new_n318_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n316_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(KEYINPUT27), .A3(new_n325_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n301_), .B1(new_n295_), .B2(new_n309_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n317_), .B1(new_n310_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n331_), .A3(KEYINPUT98), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  INV_X1    g132(.A(G155gat), .ZN(new_n334_));
  INV_X1    g133(.A(G162gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT82), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(G155gat), .A3(G162gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n333_), .B1(new_n339_), .B2(KEYINPUT1), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n336_), .A2(new_n341_), .A3(new_n338_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT83), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n336_), .A2(KEYINPUT83), .A3(new_n341_), .A4(new_n338_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n333_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT85), .B1(new_n347_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT2), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT2), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n356_), .B1(new_n347_), .B2(KEYINPUT85), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n355_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n349_), .B(KEYINPUT3), .Z(new_n359_));
  OAI211_X1 g158(.A(new_n339_), .B(new_n352_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n351_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT29), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n362_), .B(new_n363_), .C1(new_n306_), .C2(new_n305_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G78gat), .B(G106gat), .Z(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n351_), .B2(new_n360_), .ZN(new_n367_));
  OAI211_X1 g166(.A(G228gat), .B(G233gat), .C1(new_n367_), .C2(new_n302_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n364_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n365_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT92), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n364_), .A2(new_n368_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n365_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT92), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n364_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n361_), .A2(KEYINPUT29), .ZN(new_n378_));
  XOR2_X1   g177(.A(G22gat), .B(G50gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n378_), .B(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n376_), .B2(KEYINPUT91), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n371_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n371_), .B2(new_n377_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n327_), .A2(new_n332_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT99), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G127gat), .B(G134gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G120gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT81), .B(G113gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(new_n351_), .A3(new_n360_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n390_), .B(new_n391_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n361_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n395_), .A3(KEYINPUT4), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT96), .B1(new_n395_), .B2(KEYINPUT4), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n361_), .A2(new_n394_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n396_), .A2(new_n398_), .A3(new_n399_), .A4(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G57gat), .B(G85gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n393_), .A2(new_n395_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n397_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n403_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n403_), .B2(new_n410_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT30), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n304_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT31), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n394_), .B(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n419_), .B(new_n424_), .Z(new_n425_));
  INV_X1    g224(.A(KEYINPUT99), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n327_), .A2(new_n386_), .A3(new_n332_), .A4(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n388_), .A2(new_n414_), .A3(new_n425_), .A4(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n425_), .ZN(new_n429_));
  NOR4_X1   g228(.A1(new_n386_), .A2(new_n413_), .A3(new_n326_), .A4(new_n318_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n385_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n371_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n411_), .A2(KEYINPUT33), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n310_), .A2(new_n330_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n408_), .B1(new_n409_), .B2(new_n398_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n396_), .A2(new_n402_), .A3(new_n399_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n436_), .B1(new_n437_), .B2(new_n398_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n411_), .A2(KEYINPUT33), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n434_), .A2(new_n435_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n301_), .A2(KEYINPUT32), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n295_), .A2(new_n309_), .A3(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n314_), .A2(new_n315_), .ZN(new_n443_));
  OAI221_X1 g242(.A(new_n442_), .B1(new_n443_), .B2(new_n441_), .C1(new_n412_), .C2(new_n411_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n433_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n429_), .B1(new_n430_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n428_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G230gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(G57gat), .ZN(new_n449_));
  INV_X1    g248(.A(G64gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G57gat), .A2(G64gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT11), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G71gat), .B(G78gat), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT11), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n451_), .A2(new_n457_), .A3(new_n452_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n455_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT8), .ZN(new_n462_));
  INV_X1    g261(.A(G85gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n297_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n462_), .B1(new_n466_), .B2(KEYINPUT65), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT7), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G99gat), .A2(G106gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n471_), .A2(new_n474_), .A3(new_n475_), .A4(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n466_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n468_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT10), .B(G99gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT64), .B(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n474_), .A2(new_n475_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n465_), .A2(KEYINPUT9), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n464_), .A2(KEYINPUT9), .A3(new_n465_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n467_), .A2(new_n478_), .A3(new_n477_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n480_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n461_), .A2(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n460_), .A2(new_n488_), .A3(new_n480_), .A4(new_n487_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n448_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT66), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n487_), .A2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n484_), .A2(new_n486_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n495_), .A2(KEYINPUT66), .A3(new_n483_), .A4(new_n485_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n480_), .A2(new_n488_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n460_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n491_), .A2(KEYINPUT12), .ZN(new_n500_));
  AOI22_X1  g299(.A1(KEYINPUT12), .A2(new_n499_), .B1(new_n500_), .B2(new_n490_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n492_), .B1(new_n501_), .B2(new_n448_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G120gat), .B(G148gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT68), .ZN(new_n504_));
  XOR2_X1   g303(.A(G176gat), .B(G204gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT69), .B1(new_n502_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n500_), .A2(new_n490_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n494_), .A2(new_n496_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n480_), .A2(new_n488_), .ZN(new_n512_));
  OAI211_X1 g311(.A(KEYINPUT12), .B(new_n461_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n513_), .A3(new_n448_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n492_), .ZN(new_n515_));
  AND4_X1   g314(.A1(KEYINPUT69), .A2(new_n514_), .A3(new_n515_), .A4(new_n508_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n502_), .B2(new_n508_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT13), .Z(new_n519_));
  XNOR2_X1  g318(.A(G29gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G50gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT71), .B(G43gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G50gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n520_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n522_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529_));
  INV_X1    g328(.A(G1gat), .ZN(new_n530_));
  INV_X1    g329(.A(G8gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT14), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G8gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n528_), .B(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(G229gat), .A3(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n528_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n535_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n523_), .A2(new_n527_), .A3(KEYINPUT15), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n528_), .A2(new_n535_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n537_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G169gat), .B(G197gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n537_), .A2(new_n545_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n519_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n489_), .B1(new_n523_), .B2(new_n527_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT35), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n511_), .A2(new_n512_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n539_), .A2(new_n541_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n557_), .B(new_n561_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(new_n556_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n560_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n564_), .B(KEYINPUT73), .C1(new_n566_), .C2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G218gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT72), .B(G190gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT36), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n564_), .A2(KEYINPUT73), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n569_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(KEYINPUT36), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT74), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n569_), .A2(new_n580_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n578_), .A2(new_n579_), .A3(KEYINPUT37), .A4(new_n581_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n535_), .B(new_n587_), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(new_n460_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(G211gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT16), .B(G183gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n589_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n593_), .B(KEYINPUT17), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n589_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n586_), .A2(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n447_), .A2(new_n555_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n530_), .A3(new_n413_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT38), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n555_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n578_), .A2(new_n581_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI211_X1 g406(.A(new_n599_), .B(new_n607_), .C1(new_n428_), .C2(new_n446_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n414_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n603_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT101), .Z(G1324gat));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n327_), .A2(new_n332_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n605_), .A2(new_n614_), .A3(new_n608_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n616_), .A3(G8gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n615_), .B2(G8gat), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n613_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(KEYINPUT39), .A3(new_n617_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n601_), .A2(new_n531_), .A3(new_n614_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n620_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT40), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n620_), .A2(new_n622_), .A3(new_n626_), .A4(new_n623_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  OAI21_X1  g429(.A(G15gat), .B1(new_n609_), .B2(new_n429_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT41), .Z(new_n632_));
  INV_X1    g431(.A(G15gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n601_), .A2(new_n633_), .A3(new_n425_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT105), .Z(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(G1326gat));
  OAI21_X1  g435(.A(G22gat), .B1(new_n609_), .B2(new_n386_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT42), .ZN(new_n638_));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n601_), .A2(new_n639_), .A3(new_n433_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1327gat));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n447_), .B2(new_n586_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n586_), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT43), .B(new_n645_), .C1(new_n428_), .C2(new_n446_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n647_), .A2(KEYINPUT44), .A3(new_n605_), .A4(new_n599_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n605_), .B(new_n599_), .C1(new_n644_), .C2(new_n646_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n642_), .B1(new_n652_), .B2(new_n414_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n648_), .A2(new_n651_), .A3(KEYINPUT106), .A4(new_n413_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(G29gat), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n606_), .B1(new_n428_), .B2(new_n446_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n555_), .A3(new_n599_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n414_), .A2(G29gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  INV_X1    g458(.A(new_n614_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G36gat), .B1(new_n652_), .B2(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n657_), .A2(G36gat), .A3(new_n660_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT45), .Z(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(KEYINPUT46), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  NAND2_X1  g467(.A1(new_n425_), .A2(G43gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n657_), .A2(new_n429_), .ZN(new_n670_));
  OAI22_X1  g469(.A1(new_n652_), .A2(new_n669_), .B1(G43gat), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g471(.A(G50gat), .B1(new_n652_), .B2(new_n386_), .ZN(new_n673_));
  OR3_X1    g472(.A1(new_n657_), .A2(G50gat), .A3(new_n386_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1331gat));
  NAND2_X1  g474(.A1(new_n600_), .A2(new_n519_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n676_), .A2(new_n677_), .B1(new_n428_), .B2(new_n446_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n678_), .B(new_n554_), .C1(new_n677_), .C2(new_n676_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT108), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n449_), .B1(new_n680_), .B2(new_n414_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT109), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT109), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n518_), .B(KEYINPUT13), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(new_n553_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n608_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT110), .B(G57gat), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n414_), .A2(new_n687_), .ZN(new_n688_));
  AOI22_X1  g487(.A1(new_n682_), .A2(new_n683_), .B1(new_n686_), .B2(new_n688_), .ZN(G1332gat));
  AOI21_X1  g488(.A(new_n450_), .B1(new_n686_), .B2(new_n614_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT48), .Z(new_n691_));
  INV_X1    g490(.A(new_n680_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n450_), .A3(new_n614_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1333gat));
  INV_X1    g493(.A(G71gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n686_), .B2(new_n425_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT49), .Z(new_n697_));
  NAND2_X1  g496(.A1(new_n425_), .A2(new_n695_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT111), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n680_), .B2(new_n699_), .ZN(G1334gat));
  INV_X1    g499(.A(G78gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n692_), .A2(new_n701_), .A3(new_n433_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n686_), .B2(new_n433_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n703_), .A2(new_n704_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1335gat));
  NAND2_X1  g506(.A1(new_n685_), .A2(new_n599_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n644_), .A2(new_n646_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(KEYINPUT113), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(KEYINPUT113), .B2(new_n709_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n414_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n656_), .A2(new_n599_), .A3(new_n685_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n463_), .A3(new_n413_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT114), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT114), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n712_), .A2(new_n717_), .A3(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1336gat));
  AOI21_X1  g518(.A(G92gat), .B1(new_n713_), .B2(new_n614_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n711_), .A2(new_n660_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g521(.A(G99gat), .B1(new_n711_), .B2(new_n429_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n713_), .A2(new_n481_), .A3(new_n425_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT51), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(new_n727_), .A3(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1338gat));
  NOR2_X1   g528(.A1(new_n708_), .A2(new_n386_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n730_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI211_X1 g532(.A(KEYINPUT115), .B(new_n730_), .C1(new_n644_), .C2(new_n646_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(G106gat), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT52), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n733_), .A2(new_n737_), .A3(G106gat), .A4(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n713_), .A2(new_n482_), .A3(new_n433_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  INV_X1    g544(.A(KEYINPUT120), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n388_), .A2(new_n413_), .A3(new_n425_), .A4(new_n427_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n514_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(KEYINPUT117), .A2(G230gat), .A3(G233gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n501_), .A2(KEYINPUT55), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n750_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n510_), .A2(new_n513_), .A3(KEYINPUT55), .A4(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n508_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n752_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n752_), .A2(KEYINPUT56), .A3(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n553_), .B1(new_n509_), .B2(new_n516_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n553_), .B(KEYINPUT116), .C1(new_n509_), .C2(new_n516_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n536_), .A2(new_n543_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n542_), .A2(new_n544_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n769_), .B(new_n549_), .C1(new_n770_), .C2(new_n543_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(new_n552_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n518_), .A2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n761_), .A2(new_n764_), .A3(KEYINPUT118), .A4(new_n765_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n768_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n606_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(KEYINPUT119), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(KEYINPUT57), .A3(new_n606_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n761_), .A2(new_n517_), .A3(new_n772_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n781_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n586_), .A3(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n778_), .A2(new_n779_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT57), .B1(new_n775_), .B2(new_n606_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(KEYINPUT119), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n599_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n600_), .A2(new_n554_), .A3(new_n684_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT54), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n747_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT59), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n746_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n747_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n795_), .B(KEYINPUT57), .C1(new_n775_), .C2(new_n606_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n779_), .A2(new_n784_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n787_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n598_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n789_), .B(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n794_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n793_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n599_), .B1(new_n797_), .B2(new_n786_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n806_), .A2(KEYINPUT121), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(KEYINPUT121), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n790_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n805_), .A2(G113gat), .A3(new_n553_), .A4(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n803_), .B2(new_n554_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1340gat));
  NOR3_X1   g613(.A1(new_n791_), .A2(new_n746_), .A3(new_n792_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT120), .B1(new_n803_), .B2(KEYINPUT59), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n519_), .B(new_n810_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G120gat), .ZN(new_n818_));
  INV_X1    g617(.A(G120gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n684_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n791_), .B(new_n820_), .C1(KEYINPUT60), .C2(new_n819_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(G1341gat));
  NAND4_X1  g621(.A1(new_n805_), .A2(G127gat), .A3(new_n598_), .A4(new_n810_), .ZN(new_n823_));
  INV_X1    g622(.A(G127gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n803_), .B2(new_n599_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1342gat));
  NAND4_X1  g625(.A1(new_n805_), .A2(G134gat), .A3(new_n586_), .A4(new_n810_), .ZN(new_n827_));
  INV_X1    g626(.A(G134gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n803_), .B2(new_n606_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1343gat));
  NAND2_X1  g629(.A1(new_n798_), .A2(new_n799_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n802_), .B1(new_n831_), .B2(new_n599_), .ZN(new_n832_));
  NOR4_X1   g631(.A1(new_n832_), .A2(new_n425_), .A3(new_n614_), .A4(new_n386_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n413_), .A3(new_n553_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n413_), .A3(new_n519_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g636(.A1(new_n833_), .A2(new_n413_), .A3(new_n598_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(new_n334_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n838_), .B(new_n841_), .ZN(G1346gat));
  NAND3_X1  g641(.A1(new_n833_), .A2(new_n413_), .A3(new_n607_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n335_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n833_), .A2(G162gat), .A3(new_n413_), .A4(new_n586_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1347gat));
  NOR2_X1   g645(.A1(new_n660_), .A2(new_n413_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n425_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n433_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n809_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G169gat), .B1(new_n850_), .B2(new_n554_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n850_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n854_), .A2(new_n553_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT62), .B(G169gat), .C1(new_n850_), .C2(new_n554_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(new_n855_), .A3(new_n856_), .ZN(G1348gat));
  AOI21_X1  g656(.A(G176gat), .B1(new_n854_), .B2(new_n519_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n848_), .ZN(new_n859_));
  NOR4_X1   g658(.A1(new_n832_), .A2(new_n207_), .A3(new_n684_), .A4(new_n433_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(G1349gat));
  INV_X1    g660(.A(new_n270_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n790_), .A2(new_n599_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n863_), .A2(KEYINPUT123), .A3(new_n849_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT123), .B1(new_n863_), .B2(new_n849_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n862_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n213_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n809_), .A2(new_n598_), .A3(new_n867_), .A4(new_n849_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1350gat));
  NAND3_X1  g670(.A1(new_n854_), .A2(new_n212_), .A3(new_n607_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G190gat), .B1(new_n850_), .B2(new_n645_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1351gat));
  NAND2_X1  g673(.A1(new_n788_), .A2(new_n790_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n875_), .A2(new_n429_), .A3(new_n433_), .A4(new_n847_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n554_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n242_), .ZN(G1352gat));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n684_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT125), .B(G204gat), .Z(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1353gat));
  NAND2_X1  g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n598_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n876_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT126), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n884_), .B(new_n886_), .ZN(G1354gat));
  NOR2_X1   g686(.A1(new_n876_), .A2(new_n606_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(G218gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n876_), .A2(new_n645_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(G218gat), .B2(new_n890_), .ZN(G1355gat));
endmodule


