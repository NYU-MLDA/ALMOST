//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT94), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT22), .B(G169gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n210_), .B2(new_n208_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n204_), .A2(new_n205_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n209_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n207_), .A2(new_n208_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n215_), .A2(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n219_), .B(new_n203_), .C1(KEYINPUT24), .C2(new_n216_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G227gat), .A2(G233gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT96), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n225_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT95), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n223_), .B(new_n231_), .Z(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT30), .B(G15gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(G71gat), .B(G99gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT31), .B(G43gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n232_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G78gat), .B(G106gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT101), .Z(new_n240_));
  NOR2_X1   g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(KEYINPUT1), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(KEYINPUT1), .B2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G141gat), .A2(G148gat), .ZN(new_n245_));
  OR2_X1    g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n245_), .B(KEYINPUT2), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT97), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(KEYINPUT3), .ZN(new_n250_));
  OR3_X1    g049(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n241_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n242_), .A3(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n250_), .A2(new_n251_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n249_), .B1(new_n255_), .B2(new_n248_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n247_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n257_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT28), .B1(new_n257_), .B2(KEYINPUT29), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G22gat), .B(G50gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n240_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n263_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n240_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n261_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n257_), .A2(KEYINPUT29), .ZN(new_n268_));
  XOR2_X1   g067(.A(G211gat), .B(G218gat), .Z(new_n269_));
  INV_X1    g068(.A(KEYINPUT99), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT21), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G228gat), .A2(G233gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT98), .Z(new_n278_));
  OR2_X1    g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n268_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT100), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n273_), .B(KEYINPUT100), .C1(new_n272_), .C2(new_n275_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(new_n268_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n280_), .B1(new_n286_), .B2(new_n278_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n264_), .A2(new_n267_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n231_), .A2(new_n257_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n226_), .A2(new_n229_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n247_), .B(new_n296_), .C1(new_n254_), .C2(new_n256_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n294_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT4), .B1(new_n231_), .B2(new_n257_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n293_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT102), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n295_), .A2(new_n301_), .A3(new_n292_), .A4(new_n297_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G29gat), .ZN(new_n303_));
  INV_X1    g102(.A(G85gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT0), .B(G57gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n295_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT102), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n300_), .A2(new_n302_), .A3(new_n308_), .A4(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT103), .B(KEYINPUT33), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT104), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT19), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n282_), .A2(new_n283_), .A3(new_n213_), .A4(new_n220_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT20), .ZN(new_n319_));
  INV_X1    g118(.A(new_n276_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n204_), .A2(new_n211_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n220_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n317_), .B1(new_n318_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n282_), .A2(new_n283_), .B1(new_n213_), .B2(new_n220_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n320_), .B2(new_n322_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n317_), .A3(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331_));
  INV_X1    g130(.A(G92gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT18), .B(G64gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n325_), .A2(new_n330_), .A3(new_n336_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n326_), .A2(new_n328_), .A3(new_n316_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n335_), .B1(new_n338_), .B2(new_n324_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n295_), .A2(new_n293_), .A3(new_n297_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n307_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n298_), .A2(new_n299_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(new_n292_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT104), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n311_), .A2(new_n346_), .A3(new_n312_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n310_), .A2(new_n302_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n348_), .A2(KEYINPUT33), .A3(new_n308_), .A4(new_n300_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n314_), .A2(new_n345_), .A3(new_n347_), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n300_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n307_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n311_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n317_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n318_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n325_), .A2(new_n330_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n336_), .A2(KEYINPUT32), .ZN(new_n358_));
  MUX2_X1   g157(.A(new_n356_), .B(new_n357_), .S(new_n358_), .Z(new_n359_));
  NAND2_X1  g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n291_), .B1(new_n350_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n287_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n266_), .B1(new_n265_), .B2(new_n261_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n262_), .A2(new_n240_), .A3(new_n263_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n365_), .A2(new_n352_), .A3(new_n311_), .A4(new_n288_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n335_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT105), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(new_n367_), .B2(new_n337_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT27), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n340_), .A2(KEYINPUT27), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n366_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n238_), .B1(new_n361_), .B2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n238_), .A2(new_n291_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n353_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(new_n374_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G1gat), .B(G8gat), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(G15gat), .A2(G22gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G15gat), .A2(G22gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT14), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(G1gat), .B2(G8gat), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n387_), .A2(new_n389_), .A3(KEYINPUT84), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G15gat), .B(G22gat), .ZN(new_n392_));
  INV_X1    g191(.A(G1gat), .ZN(new_n393_));
  INV_X1    g192(.A(G8gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT14), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n384_), .B1(new_n390_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT84), .B1(new_n387_), .B2(new_n389_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n392_), .A2(new_n391_), .A3(new_n395_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n383_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G231gat), .A2(G233gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n404_));
  XOR2_X1   g203(.A(G183gat), .B(G211gat), .Z(new_n405_));
  XNOR2_X1  g204(.A(G127gat), .B(G155gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n404_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n403_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G71gat), .B(G78gat), .ZN(new_n413_));
  INV_X1    g212(.A(G57gat), .ZN(new_n414_));
  INV_X1    g213(.A(G64gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G57gat), .A2(G64gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT70), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT70), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n420_), .A3(new_n417_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n413_), .B1(new_n422_), .B2(KEYINPUT11), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT11), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n419_), .A2(new_n424_), .A3(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(KEYINPUT11), .A3(new_n413_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n412_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n409_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n430_), .B1(KEYINPUT17), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n412_), .A2(new_n429_), .ZN(new_n433_));
  OR3_X1    g232(.A1(new_n432_), .A2(KEYINPUT87), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT87), .B1(new_n432_), .B2(new_n433_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G190gat), .B(G218gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G134gat), .B(G162gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n440_), .A2(KEYINPUT36), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(KEYINPUT36), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n445_));
  NAND2_X1  g244(.A1(G232gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(KEYINPUT76), .B(KEYINPUT35), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G85gat), .B(G92gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT68), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n304_), .A2(G92gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n332_), .A2(G85gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT68), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT8), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT65), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT6), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G99gat), .A2(G106gat), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n461_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n464_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n459_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n464_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n462_), .A2(KEYINPUT6), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n460_), .A2(KEYINPUT65), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n461_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT66), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT67), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT7), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT67), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  AOI211_X1 g279(.A(G99gat), .B(G106gat), .C1(new_n476_), .C2(KEYINPUT7), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n458_), .B1(new_n474_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n465_), .A2(new_n466_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n477_), .A2(new_n475_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n475_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n456_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT69), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n457_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(KEYINPUT69), .B(new_n456_), .C1(new_n484_), .C2(new_n487_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n483_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT9), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT10), .B(G99gat), .ZN(new_n494_));
  OAI22_X1  g293(.A1(new_n493_), .A2(new_n450_), .B1(new_n494_), .B2(G106gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT64), .B(G85gat), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n496_), .A2(KEYINPUT9), .A3(new_n332_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n474_), .A2(KEYINPUT71), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT71), .B1(new_n474_), .B2(new_n498_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n492_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT77), .ZN(new_n503_));
  INV_X1    g302(.A(G50gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G43gat), .ZN(new_n505_));
  INV_X1    g304(.A(G43gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G50gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n507_), .A3(new_n503_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G29gat), .B(G36gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n511_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n505_), .A2(new_n507_), .A3(new_n503_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(new_n508_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n512_), .A2(new_n515_), .A3(KEYINPUT15), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT15), .B1(new_n512_), .B2(new_n515_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT78), .B1(new_n502_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n500_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n474_), .A2(KEYINPUT71), .A3(new_n498_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n465_), .A2(new_n466_), .A3(new_n459_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT66), .B1(new_n471_), .B2(new_n472_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n482_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n458_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n471_), .A2(new_n472_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n528_), .A2(new_n482_), .B1(new_n455_), .B2(new_n452_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT8), .B1(new_n529_), .B2(KEYINPUT69), .ZN(new_n530_));
  INV_X1    g329(.A(new_n491_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n527_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n522_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT78), .ZN(new_n534_));
  INV_X1    g333(.A(new_n518_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n519_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n512_), .A2(new_n515_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n474_), .A2(new_n498_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT79), .ZN(new_n542_));
  INV_X1    g341(.A(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n488_), .A2(new_n489_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(KEYINPUT8), .A3(new_n491_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n545_), .B2(new_n527_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT79), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n539_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n542_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n447_), .A2(new_n448_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AND4_X1   g350(.A1(new_n449_), .A2(new_n537_), .A3(new_n549_), .A4(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n519_), .B2(new_n536_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n449_), .B1(new_n553_), .B2(new_n549_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n444_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n519_), .A2(new_n536_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n549_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n448_), .B(new_n447_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n553_), .A2(new_n449_), .A3(new_n549_), .ZN(new_n559_));
  XOR2_X1   g358(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n441_), .B(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n443_), .B(KEYINPUT82), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n565_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n563_), .B1(new_n566_), .B2(new_n562_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n564_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AOI211_X1 g368(.A(KEYINPUT83), .B(new_n563_), .C1(new_n566_), .C2(new_n562_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n436_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n398_), .A2(new_n383_), .A3(new_n399_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n383_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n538_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n397_), .A2(new_n400_), .A3(new_n512_), .A4(new_n515_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(KEYINPUT88), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT88), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n401_), .A2(new_n579_), .A3(new_n538_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n576_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n401_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n577_), .B(KEYINPUT89), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n575_), .A3(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n581_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT93), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n581_), .A2(new_n585_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT90), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n581_), .A2(KEYINPUT90), .A3(new_n585_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n588_), .B(KEYINPUT91), .Z(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT92), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n581_), .A2(KEYINPUT90), .A3(new_n585_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT90), .B1(new_n581_), .B2(new_n585_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT92), .B(new_n597_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n591_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n546_), .B2(new_n428_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G230gat), .A2(G233gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n532_), .A2(new_n428_), .A3(new_n540_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n428_), .A2(new_n604_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n492_), .B2(new_n501_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n606_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n607_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n428_), .B1(new_n532_), .B2(new_n540_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n611_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(G204gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT73), .B(G176gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n610_), .A2(new_n614_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT74), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT74), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n610_), .A2(new_n614_), .A3(new_n623_), .A4(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n610_), .A2(new_n614_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n620_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(KEYINPUT13), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(KEYINPUT13), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n603_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n382_), .A2(new_n571_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(G1gat), .A3(new_n378_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n635_), .A2(KEYINPUT38), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(KEYINPUT38), .ZN(new_n637_));
  INV_X1    g436(.A(new_n436_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n555_), .A2(new_n562_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n381_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n632_), .B(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n645_), .B2(new_n378_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n636_), .A2(new_n637_), .A3(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(new_n379_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n633_), .A2(new_n394_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  INV_X1    g449(.A(new_n645_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n648_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n650_), .B1(new_n652_), .B2(G8gat), .ZN(new_n653_));
  AOI211_X1 g452(.A(KEYINPUT39), .B(new_n394_), .C1(new_n651_), .C2(new_n648_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n649_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(G1325gat));
  OAI21_X1  g456(.A(G15gat), .B1(new_n645_), .B2(new_n238_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(KEYINPUT41), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(KEYINPUT41), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n634_), .A2(G15gat), .A3(new_n238_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n659_), .A2(new_n660_), .A3(new_n661_), .ZN(G1326gat));
  INV_X1    g461(.A(new_n291_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G22gat), .B1(new_n645_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n663_), .A2(G22gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n634_), .B2(new_n666_), .ZN(G1327gat));
  NOR2_X1   g466(.A1(new_n569_), .A2(new_n570_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n381_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n381_), .A2(KEYINPUT43), .A3(new_n668_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n638_), .A4(new_n644_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n436_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n676_), .A2(KEYINPUT44), .A3(new_n644_), .A4(new_n672_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n677_), .A3(new_n353_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G29gat), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n382_), .A2(new_n632_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n436_), .A2(new_n639_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT107), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n378_), .A2(G29gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n679_), .B1(new_n683_), .B2(new_n684_), .ZN(G1328gat));
  NAND3_X1  g484(.A1(new_n675_), .A2(new_n677_), .A3(new_n648_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G36gat), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n379_), .A2(G36gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n680_), .A2(new_n682_), .A3(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT45), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n687_), .B(new_n690_), .C1(KEYINPUT108), .C2(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1329gat));
  NOR2_X1   g494(.A1(new_n238_), .A2(new_n506_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n675_), .A2(new_n677_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT109), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n675_), .A2(new_n677_), .A3(new_n699_), .A4(new_n696_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n506_), .B1(new_n683_), .B2(new_n238_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT47), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n698_), .A2(new_n704_), .A3(new_n700_), .A4(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1330gat));
  NAND3_X1  g505(.A1(new_n675_), .A2(new_n677_), .A3(new_n291_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G50gat), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n680_), .A2(new_n504_), .A3(new_n291_), .A4(new_n682_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT110), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n630_), .A2(new_n631_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n603_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(new_n381_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(new_n641_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(G57gat), .A3(new_n353_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n566_), .A2(new_n562_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT37), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT83), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n567_), .A2(new_n568_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n564_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n718_), .A2(new_n436_), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n414_), .B1(new_n728_), .B2(new_n378_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n720_), .A2(new_n721_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n722_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT112), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n722_), .A2(new_n733_), .A3(new_n729_), .A4(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1332gat));
  AOI21_X1  g534(.A(new_n415_), .B1(new_n719_), .B2(new_n648_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n648_), .A2(new_n415_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n728_), .B2(new_n739_), .ZN(G1333gat));
  INV_X1    g539(.A(new_n719_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G71gat), .B1(new_n741_), .B2(new_n238_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT49), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n238_), .A2(G71gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n728_), .B2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n741_), .B2(new_n663_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT50), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n663_), .A2(G78gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n728_), .B2(new_n748_), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n718_), .A2(new_n682_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n353_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n676_), .A2(new_n672_), .A3(new_n717_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n753_), .A2(new_n496_), .A3(new_n378_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1336gat));
  OAI21_X1  g554(.A(new_n332_), .B1(new_n750_), .B2(new_n379_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n648_), .A2(G92gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n753_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT114), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n753_), .B2(new_n238_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n238_), .A2(new_n494_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n750_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n762_), .B(new_n763_), .Z(G1338gat));
  OR3_X1    g563(.A1(new_n750_), .A2(G106gat), .A3(new_n663_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n676_), .A2(new_n291_), .A3(new_n672_), .A4(new_n717_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n765_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n625_), .A2(new_n603_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n533_), .A2(new_n608_), .B1(new_n546_), .B2(new_n428_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n606_), .B1(new_n776_), .B2(new_n605_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n610_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n776_), .A2(KEYINPUT55), .A3(new_n606_), .A4(new_n605_), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n775_), .B(new_n620_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n774_), .B1(new_n781_), .B2(KEYINPUT116), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n607_), .B(new_n609_), .C1(new_n613_), .C2(KEYINPUT12), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n778_), .B1(new_n783_), .B2(new_n611_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n610_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n780_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n627_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n775_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT56), .B(new_n627_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n782_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n576_), .A2(new_n584_), .A3(new_n580_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n582_), .A2(new_n575_), .A3(new_n583_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n588_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n591_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n640_), .B1(new_n793_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n773_), .B1(new_n801_), .B2(KEYINPUT57), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n799_), .B1(new_n782_), .B2(new_n792_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT117), .B(new_n803_), .C1(new_n804_), .C2(new_n640_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n597_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT92), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n601_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n591_), .A2(new_n809_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n791_), .B2(new_n790_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n779_), .A2(new_n780_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n627_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n781_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n811_), .B1(new_n814_), .B2(new_n790_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n639_), .C1(new_n815_), .C2(new_n799_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n569_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n798_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n813_), .B2(new_n781_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT58), .B(new_n818_), .C1(new_n813_), .C2(new_n781_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n817_), .A2(new_n821_), .A3(new_n726_), .A4(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n802_), .A2(new_n805_), .A3(new_n816_), .A4(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n638_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n603_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT54), .B1(new_n571_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n631_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n629_), .A2(KEYINPUT13), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n603_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n727_), .A2(new_n831_), .A3(new_n832_), .A4(new_n436_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n828_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n825_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n648_), .A2(new_n378_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n377_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT59), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n803_), .B1(new_n804_), .B2(new_n640_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(new_n816_), .A3(new_n823_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n638_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n834_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT59), .B1(new_n837_), .B2(KEYINPUT118), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n844_), .B(new_n845_), .C1(KEYINPUT118), .C2(new_n837_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n826_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n840_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n839_), .B2(new_n826_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1340gat));
  AND2_X1   g650(.A1(new_n828_), .A2(new_n833_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n824_), .B2(new_n638_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n837_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n715_), .B(new_n846_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G120gat), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT60), .ZN(new_n858_));
  AOI21_X1  g657(.A(G120gat), .B1(new_n715_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n860_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n858_), .B2(G120gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n854_), .A2(new_n861_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n857_), .A2(new_n864_), .ZN(G1341gat));
  NOR2_X1   g664(.A1(new_n638_), .A2(KEYINPUT120), .ZN(new_n866_));
  MUX2_X1   g665(.A(KEYINPUT120), .B(new_n866_), .S(G127gat), .Z(new_n867_));
  NAND3_X1  g666(.A1(new_n840_), .A2(new_n846_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(G127gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n839_), .B2(new_n638_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1342gat));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT121), .B(new_n872_), .C1(new_n839_), .C2(new_n639_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n853_), .A2(new_n639_), .A3(new_n837_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(G134gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT122), .B(G134gat), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n727_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n846_), .B(new_n878_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n873_), .A2(new_n876_), .A3(new_n879_), .ZN(G1343gat));
  INV_X1    g679(.A(new_n238_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n853_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n836_), .A2(new_n291_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(new_n603_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g685(.A1(new_n882_), .A2(new_n715_), .A3(new_n884_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g687(.A1(new_n882_), .A2(new_n436_), .A3(new_n884_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1346gat));
  NOR4_X1   g690(.A1(new_n853_), .A2(new_n639_), .A3(new_n881_), .A4(new_n883_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT123), .B1(new_n892_), .B2(G162gat), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n835_), .A2(new_n640_), .A3(new_n238_), .A4(new_n884_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895_));
  INV_X1    g694(.A(G162gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n882_), .A2(G162gat), .A3(new_n668_), .A4(new_n884_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n893_), .A2(new_n897_), .A3(new_n898_), .ZN(G1347gat));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n648_), .A2(new_n378_), .A3(new_n377_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n843_), .B2(new_n834_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(new_n210_), .A3(new_n603_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n207_), .B1(new_n902_), .B2(new_n603_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(KEYINPUT62), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n826_), .B(new_n901_), .C1(new_n843_), .C2(new_n834_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n207_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n900_), .B1(new_n905_), .B2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n904_), .A2(KEYINPUT62), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n907_), .B1(new_n906_), .B2(new_n207_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(KEYINPUT124), .A4(new_n903_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(G1348gat));
  AOI21_X1  g712(.A(G176gat), .B1(new_n902_), .B2(new_n715_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n853_), .A2(new_n901_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n716_), .A2(new_n208_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1349gat));
  AOI21_X1  g716(.A(G183gat), .B1(new_n915_), .B2(new_n436_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n901_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n844_), .A2(new_n919_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n920_), .A2(new_n638_), .A3(new_n217_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n918_), .A2(new_n921_), .ZN(G1350gat));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n727_), .ZN(new_n923_));
  INV_X1    g722(.A(G190gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n640_), .A2(new_n218_), .ZN(new_n925_));
  OAI22_X1  g724(.A1(new_n923_), .A2(new_n924_), .B1(new_n920_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  OAI221_X1 g727(.A(new_n928_), .B1(new_n920_), .B2(new_n925_), .C1(new_n923_), .C2(new_n924_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1351gat));
  NOR2_X1   g729(.A1(new_n379_), .A2(new_n366_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n882_), .A2(new_n603_), .A3(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G197gat), .ZN(G1352gat));
  NOR4_X1   g732(.A1(new_n853_), .A2(new_n366_), .A3(new_n379_), .A4(new_n881_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n715_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(G204gat), .ZN(new_n936_));
  INV_X1    g735(.A(G204gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n934_), .A2(new_n937_), .A3(new_n715_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1353gat));
  XNOR2_X1  g738(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n940_), .B(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n638_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n943_));
  AND3_X1   g742(.A1(new_n934_), .A2(new_n942_), .A3(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n942_), .B1(new_n934_), .B2(new_n943_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1354gat));
  AOI21_X1  g745(.A(G218gat), .B1(new_n934_), .B2(new_n640_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n668_), .A2(G218gat), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n934_), .B2(new_n948_), .ZN(G1355gat));
endmodule


