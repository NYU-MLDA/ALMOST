//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_;
  INV_X1    g000(.A(G233gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n202_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(G204gat), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  INV_X1    g009(.A(G204gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G197gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n211_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n210_), .B1(G197gat), .B2(G204gat), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n215_), .A2(KEYINPUT86), .A3(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT86), .B1(new_n215_), .B2(new_n216_), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n213_), .B(new_n214_), .C1(new_n217_), .C2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n212_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT85), .B(G197gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(G204gat), .ZN(new_n222_));
  OR3_X1    g021(.A1(new_n222_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT89), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT82), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT1), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n227_), .B(new_n228_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n228_), .B(KEYINPUT2), .Z(new_n234_));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n226_), .B(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n231_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n233_), .B1(new_n237_), .B2(new_n230_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT29), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n206_), .B1(new_n225_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT90), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n243_), .B(new_n206_), .C1(new_n225_), .C2(new_n240_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n213_), .A2(new_n214_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n218_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n215_), .A2(KEYINPUT86), .A3(new_n216_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n222_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT87), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT87), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n219_), .A2(new_n223_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n206_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(new_n239_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT88), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT88), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n254_), .A2(new_n258_), .A3(new_n255_), .A4(new_n239_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n245_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G78gat), .B(G106gat), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n238_), .A2(KEYINPUT29), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT83), .B(KEYINPUT28), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G22gat), .B(G50gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n265_), .B(new_n268_), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT91), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n260_), .A2(new_n242_), .A3(new_n244_), .A4(new_n262_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n264_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n262_), .B1(new_n245_), .B2(new_n260_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n272_), .A2(new_n269_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n270_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT20), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT77), .ZN(new_n279_));
  INV_X1    g078(.A(G190gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(KEYINPUT26), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT25), .B(G183gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(G190gat), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n281_), .B(new_n282_), .C1(new_n283_), .C2(new_n279_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT78), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT23), .ZN(new_n287_));
  OR3_X1    g086(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n288_));
  OR2_X1    g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(KEYINPUT24), .A3(new_n290_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n287_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n280_), .A2(KEYINPUT26), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(G190gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT77), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n281_), .A4(new_n282_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n285_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT79), .B(G176gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT22), .B(G169gat), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n300_), .A2(new_n301_), .B1(G169gat), .B2(G176gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT80), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(new_n286_), .B2(KEYINPUT23), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n287_), .B2(new_n303_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n302_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n299_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n278_), .B1(new_n254_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n224_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n291_), .A2(new_n288_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n283_), .A2(new_n282_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n286_), .B(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(KEYINPUT80), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n314_), .B(new_n315_), .C1(new_n318_), .C2(new_n304_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n300_), .A2(new_n301_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n290_), .B(KEYINPUT93), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n320_), .B(new_n321_), .C1(new_n317_), .C2(new_n306_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n312_), .B1(new_n313_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n309_), .A2(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n299_), .A2(new_n307_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n251_), .A2(new_n326_), .A3(new_n253_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n319_), .A2(new_n322_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n278_), .B1(new_n224_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT94), .B1(new_n330_), .B2(new_n312_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT94), .ZN(new_n332_));
  INV_X1    g131(.A(new_n312_), .ZN(new_n333_));
  AOI211_X1 g132(.A(new_n332_), .B(new_n333_), .C1(new_n327_), .C2(new_n329_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n325_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G8gat), .B(G36gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G92gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT18), .B(G64gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n325_), .B(new_n339_), .C1(new_n331_), .C2(new_n334_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT27), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n327_), .A2(new_n329_), .A3(new_n333_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT97), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n327_), .A2(KEYINPUT97), .A3(new_n329_), .A4(new_n333_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT96), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n328_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n323_), .A2(KEYINPUT96), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n224_), .A2(KEYINPUT89), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n224_), .A2(KEYINPUT89), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n350_), .B(new_n351_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n333_), .B1(new_n309_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n340_), .B1(new_n348_), .B2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n356_), .A2(KEYINPUT27), .A3(new_n342_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT98), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n343_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT27), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n219_), .A2(new_n223_), .A3(new_n252_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n252_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n361_), .A2(new_n362_), .A3(new_n308_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT20), .B1(new_n313_), .B2(new_n323_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n312_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n332_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n330_), .A2(KEYINPUT94), .A3(new_n312_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n339_), .B1(new_n368_), .B2(new_n325_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n342_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n360_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n356_), .A2(KEYINPUT27), .A3(new_n342_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT98), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n277_), .B1(new_n359_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT99), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377_));
  XOR2_X1   g176(.A(G113gat), .B(G120gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n238_), .A2(new_n377_), .A3(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n238_), .B(new_n380_), .Z(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(KEYINPUT4), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n384_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  INV_X1    g188(.A(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n393_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n386_), .A2(new_n387_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n380_), .B(KEYINPUT31), .Z(new_n399_));
  XNOR2_X1  g198(.A(new_n308_), .B(KEYINPUT30), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G43gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(G15gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n401_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n399_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n409_), .B1(new_n408_), .B2(new_n407_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n407_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(KEYINPUT81), .A3(new_n399_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n277_), .B(KEYINPUT99), .C1(new_n359_), .C2(new_n373_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n376_), .A2(new_n398_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n396_), .B(KEYINPUT33), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n383_), .A2(new_n384_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n418_), .A2(KEYINPUT95), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(KEYINPUT95), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n382_), .A2(new_n385_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n419_), .A2(new_n393_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n417_), .A2(new_n422_), .A3(new_n342_), .A4(new_n341_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n339_), .A2(KEYINPUT32), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n348_), .B2(new_n355_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n397_), .B(new_n425_), .C1(new_n335_), .C2(new_n424_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n277_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n343_), .A2(new_n357_), .A3(new_n397_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n427_), .B(new_n413_), .C1(new_n277_), .C2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n416_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G99gat), .A2(G106gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT6), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n433_));
  OR3_X1    g232(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G85gat), .B(G92gat), .Z(new_n436_));
  NAND2_X1  g235(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(KEYINPUT9), .ZN(new_n441_));
  XOR2_X1   g240(.A(KEYINPUT10), .B(G99gat), .Z(new_n442_));
  INV_X1    g241(.A(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G92gat), .ZN(new_n445_));
  OR3_X1    g244(.A1(new_n390_), .A2(new_n445_), .A3(KEYINPUT9), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n441_), .A2(new_n444_), .A3(new_n446_), .A4(new_n432_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n439_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .A4(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n440_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT66), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n440_), .A2(new_n452_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G57gat), .B(G64gat), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n455_), .A2(KEYINPUT11), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(KEYINPUT11), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G71gat), .B(G78gat), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n459_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n454_), .A2(KEYINPUT12), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G230gat), .A2(G233gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT64), .Z(new_n463_));
  XOR2_X1   g262(.A(KEYINPUT67), .B(KEYINPUT12), .Z(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n450_), .B2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n450_), .A2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n450_), .B(new_n460_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n463_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G120gat), .B(G148gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G204gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT5), .B(G176gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n472_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT13), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n479_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483_));
  INV_X1    g282(.A(G36gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT68), .B(G29gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n483_), .B(G36gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n486_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492_));
  INV_X1    g291(.A(G1gat), .ZN(new_n493_));
  INV_X1    g292(.A(G8gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G1gat), .B(G8gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT75), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n487_), .A2(new_n490_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n491_), .B(KEYINPUT15), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT76), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n502_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n501_), .A2(KEYINPUT15), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n491_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n502_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT76), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n510_), .A2(new_n515_), .A3(new_n500_), .A4(new_n505_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n507_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G169gat), .B(G197gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n507_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n482_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n430_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT72), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT34), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n454_), .A2(new_n508_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n491_), .A2(new_n440_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT69), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n532_), .A2(new_n529_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT70), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n538_), .A2(KEYINPUT70), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n537_), .A2(new_n542_), .A3(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n533_), .A2(KEYINPUT70), .A3(new_n538_), .A4(new_n536_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n528_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(G162gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT71), .B(G134gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT36), .B1(new_n547_), .B2(new_n552_), .ZN(new_n553_));
  AOI211_X1 g352(.A(new_n541_), .B(new_n543_), .C1(new_n533_), .C2(new_n536_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n546_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT72), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n551_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n552_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n553_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT37), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT37), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n553_), .A2(new_n558_), .A3(new_n562_), .A4(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n460_), .B(new_n502_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT73), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n565_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G211gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT16), .B(G183gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(KEYINPUT74), .A3(KEYINPUT17), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(KEYINPUT17), .B2(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n568_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n564_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n527_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n493_), .A3(new_n397_), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n560_), .A2(KEYINPUT101), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n560_), .A2(KEYINPUT101), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(new_n579_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n527_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n589_), .A2(new_n397_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n584_), .B1(new_n493_), .B2(new_n590_), .ZN(G1324gat));
  NOR2_X1   g390(.A1(new_n359_), .A2(new_n373_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n494_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT39), .Z(new_n594_));
  NAND3_X1  g393(.A1(new_n581_), .A2(new_n494_), .A3(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g396(.A(new_n403_), .B1(new_n589_), .B2(new_n414_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT41), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n581_), .A2(new_n403_), .A3(new_n414_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(G1326gat));
  INV_X1    g400(.A(G22gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n277_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n589_), .B2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT42), .Z(new_n605_));
  NAND3_X1  g404(.A1(new_n581_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1327gat));
  INV_X1    g406(.A(new_n587_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(new_n578_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n527_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(G29gat), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n397_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n430_), .A2(new_n614_), .A3(new_n564_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n430_), .A2(new_n564_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT43), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n430_), .A2(KEYINPUT102), .A3(new_n614_), .A4(new_n564_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n526_), .A3(new_n579_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT44), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n621_), .A2(KEYINPUT44), .A3(new_n526_), .A4(new_n579_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n397_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n613_), .B1(new_n627_), .B2(G29gat), .ZN(new_n628_));
  AOI211_X1 g427(.A(KEYINPUT103), .B(new_n611_), .C1(new_n626_), .C2(new_n397_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n612_), .B1(new_n628_), .B2(new_n629_), .ZN(G1328gat));
  NOR2_X1   g429(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT46), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n624_), .A2(new_n592_), .A3(new_n625_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(G36gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n592_), .B(KEYINPUT104), .Z(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n610_), .A2(new_n484_), .A3(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT45), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n631_), .B(new_n634_), .C1(new_n636_), .C2(new_n640_), .ZN(new_n641_));
  AND4_X1   g440(.A1(new_n632_), .A2(new_n636_), .A3(new_n633_), .A4(new_n640_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1329gat));
  NAND3_X1  g442(.A1(new_n626_), .A2(G43gat), .A3(new_n414_), .ZN(new_n644_));
  INV_X1    g443(.A(G43gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n610_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(new_n413_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n644_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n644_), .B2(new_n647_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1330gat));
  NAND2_X1  g450(.A1(new_n626_), .A2(new_n603_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT107), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n626_), .A2(new_n654_), .A3(new_n603_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(G50gat), .A3(new_n655_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n277_), .A2(G50gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n646_), .B2(new_n657_), .ZN(G1331gat));
  INV_X1    g457(.A(new_n482_), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n524_), .B(new_n659_), .C1(new_n416_), .C2(new_n429_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(new_n588_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n397_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n660_), .A2(new_n580_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n398_), .A2(G57gat), .ZN(new_n664_));
  AOI22_X1  g463(.A1(new_n662_), .A2(G57gat), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT108), .Z(G1332gat));
  INV_X1    g465(.A(G64gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n661_), .B2(new_n638_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT48), .Z(new_n669_));
  NAND3_X1  g468(.A1(new_n663_), .A2(new_n667_), .A3(new_n638_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1333gat));
  INV_X1    g470(.A(G71gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n661_), .B2(new_n414_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT49), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n663_), .A2(new_n672_), .A3(new_n414_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT109), .ZN(G1334gat));
  INV_X1    g476(.A(G78gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n661_), .B2(new_n603_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT50), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n663_), .A2(new_n678_), .A3(new_n603_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1335gat));
  AND2_X1   g481(.A1(new_n660_), .A2(new_n609_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G85gat), .B1(new_n683_), .B2(new_n397_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n659_), .A2(new_n524_), .A3(new_n578_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n621_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n398_), .A2(new_n390_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(G1336gat));
  AOI21_X1  g487(.A(G92gat), .B1(new_n683_), .B2(new_n592_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n637_), .A2(new_n445_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n686_), .B2(new_n690_), .ZN(G1337gat));
  NAND2_X1  g490(.A1(new_n686_), .A2(new_n414_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n414_), .A2(new_n442_), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n692_), .A2(G99gat), .B1(new_n683_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT51), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(KEYINPUT110), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(KEYINPUT110), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1338gat));
  NAND3_X1  g497(.A1(new_n621_), .A2(new_n603_), .A3(new_n685_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n621_), .A2(KEYINPUT111), .A3(new_n603_), .A4(new_n685_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(G106gat), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT52), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT52), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n701_), .A2(new_n705_), .A3(G106gat), .A4(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n683_), .A2(new_n443_), .A3(new_n603_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT53), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT53), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n707_), .A2(new_n711_), .A3(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1339gat));
  NAND3_X1  g512(.A1(new_n580_), .A2(new_n525_), .A3(new_n659_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT54), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT116), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT58), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n461_), .A2(new_n467_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n470_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(KEYINPUT55), .A3(new_n468_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n468_), .A2(KEYINPUT55), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n476_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT56), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n721_), .A2(new_n722_), .A3(KEYINPUT56), .A4(new_n476_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n472_), .A2(new_n477_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n504_), .A2(new_n505_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n510_), .A2(new_n515_), .A3(new_n500_), .A4(new_n506_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n520_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n523_), .A2(new_n732_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n729_), .B(new_n733_), .C1(new_n727_), .C2(new_n726_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n718_), .B1(new_n728_), .B2(new_n734_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n564_), .A2(new_n735_), .A3(KEYINPUT114), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT114), .B1(new_n564_), .B2(new_n735_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n733_), .A2(new_n729_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n727_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(KEYINPUT113), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(KEYINPUT58), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n740_), .A2(new_n741_), .A3(KEYINPUT115), .A4(KEYINPUT58), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n736_), .A2(new_n737_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n478_), .A2(new_n733_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n725_), .A2(new_n727_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n524_), .A2(new_n729_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n585_), .A2(new_n751_), .A3(new_n586_), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT112), .B(KEYINPUT57), .Z(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n717_), .B1(new_n747_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT57), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n752_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n564_), .A2(new_n735_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n744_), .A2(new_n745_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n564_), .A2(new_n735_), .A3(KEYINPUT114), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT116), .A3(new_n754_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n756_), .A2(new_n759_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n716_), .B1(new_n767_), .B2(new_n579_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n376_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n397_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(KEYINPUT59), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT117), .B1(new_n768_), .B2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n765_), .A2(new_n759_), .A3(new_n754_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n579_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(new_n715_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT59), .B1(new_n776_), .B2(new_n770_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n765_), .A2(new_n754_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n758_), .B1(new_n779_), .B2(new_n717_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n578_), .B1(new_n780_), .B2(new_n766_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n778_), .B(new_n771_), .C1(new_n781_), .C2(new_n716_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n773_), .A2(new_n777_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(G113gat), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(new_n525_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n776_), .A2(new_n770_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G113gat), .B1(new_n786_), .B2(new_n524_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1340gat));
  INV_X1    g587(.A(KEYINPUT60), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n659_), .B2(G120gat), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n786_), .B(new_n790_), .C1(new_n789_), .C2(G120gat), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT118), .ZN(new_n792_));
  OAI21_X1  g591(.A(G120gat), .B1(new_n783_), .B2(new_n659_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1341gat));
  INV_X1    g593(.A(G127gat), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n783_), .A2(new_n795_), .A3(new_n579_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G127gat), .B1(new_n786_), .B2(new_n578_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1342gat));
  NAND4_X1  g597(.A1(new_n773_), .A2(new_n782_), .A3(new_n564_), .A4(new_n777_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G134gat), .ZN(new_n800_));
  INV_X1    g599(.A(G134gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n786_), .A2(new_n801_), .A3(new_n587_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n800_), .A2(KEYINPUT119), .A3(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(G1343gat));
  NOR3_X1   g606(.A1(new_n776_), .A2(new_n414_), .A3(new_n277_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n397_), .A3(new_n637_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n525_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT120), .B(G141gat), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(G1344gat));
  NOR2_X1   g611(.A1(new_n809_), .A2(new_n659_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g613(.A1(new_n809_), .A2(new_n579_), .ZN(new_n815_));
  XOR2_X1   g614(.A(KEYINPUT61), .B(G155gat), .Z(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(G1346gat));
  INV_X1    g616(.A(new_n564_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G162gat), .B1(new_n809_), .B2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n608_), .A2(G162gat), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n808_), .A2(new_n397_), .A3(new_n637_), .A4(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT121), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n819_), .A2(new_n824_), .A3(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1347gat));
  INV_X1    g625(.A(new_n768_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n637_), .A2(new_n397_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n414_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT122), .Z(new_n830_));
  NAND4_X1  g629(.A1(new_n827_), .A2(new_n524_), .A3(new_n277_), .A4(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT62), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(G169gat), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n831_), .B2(G169gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n827_), .A2(new_n277_), .A3(new_n830_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n524_), .A2(new_n301_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT123), .ZN(new_n838_));
  OAI22_X1  g637(.A1(new_n834_), .A2(new_n835_), .B1(new_n836_), .B2(new_n838_), .ZN(G1348gat));
  NOR2_X1   g638(.A1(new_n776_), .A2(new_n603_), .ZN(new_n840_));
  AND4_X1   g639(.A1(G176gat), .A2(new_n840_), .A3(new_n482_), .A4(new_n830_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n300_), .B1(new_n836_), .B2(new_n659_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n842_), .A2(KEYINPUT124), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(KEYINPUT124), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(G1349gat));
  NOR3_X1   g644(.A1(new_n836_), .A2(new_n282_), .A3(new_n579_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n830_), .A2(new_n578_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G183gat), .B1(new_n847_), .B2(new_n840_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1350gat));
  NAND4_X1  g648(.A1(new_n827_), .A2(new_n277_), .A3(new_n564_), .A4(new_n830_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT125), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(G190gat), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n850_), .B2(G190gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n587_), .A2(new_n283_), .ZN(new_n855_));
  OAI22_X1  g654(.A1(new_n853_), .A2(new_n854_), .B1(new_n836_), .B2(new_n855_), .ZN(G1351gat));
  AND2_X1   g655(.A1(new_n808_), .A2(new_n828_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n524_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n482_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n211_), .A2(KEYINPUT126), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1353gat));
  AOI21_X1  g661(.A(new_n579_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT127), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n863_), .A2(KEYINPUT127), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n857_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n866_), .B(new_n867_), .Z(G1354gat));
  AOI21_X1  g667(.A(G218gat), .B1(new_n857_), .B2(new_n587_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n564_), .A2(G218gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n857_), .B2(new_n870_), .ZN(G1355gat));
endmodule


