//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_;
  XNOR2_X1  g000(.A(KEYINPUT73), .B(G43gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G50gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G29gat), .B(G36gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G50gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n202_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n204_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n209_), .A3(KEYINPUT15), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n205_), .A2(new_n209_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NOR3_X1   g015(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n214_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT6), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT66), .A3(new_n215_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n218_), .A2(new_n220_), .A3(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G85gat), .B(G92gat), .Z(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n225_), .A2(KEYINPUT67), .A3(new_n226_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(KEYINPUT8), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT68), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n229_), .A2(new_n233_), .A3(KEYINPUT8), .A4(new_n230_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n220_), .A2(new_n215_), .A3(new_n223_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n226_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT9), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n226_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT10), .B(G99gat), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(G106gat), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n242_), .A2(new_n243_), .A3(G85gat), .A4(G92gat), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .A4(new_n220_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n240_), .A2(new_n241_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n241_), .B1(new_n240_), .B2(new_n250_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n210_), .B(new_n213_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G232gat), .A2(G233gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n254_), .B(KEYINPUT72), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT34), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n256_), .A2(KEYINPUT35), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n240_), .A2(new_n211_), .A3(new_n250_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(KEYINPUT35), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n260_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G190gat), .B(G218gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G134gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(G162gat), .Z(new_n266_));
  INV_X1    g065(.A(KEYINPUT36), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n266_), .B(new_n267_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n261_), .A2(new_n262_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT37), .B1(new_n269_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n263_), .A2(new_n268_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT37), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n271_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G57gat), .B(G64gat), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT11), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT11), .ZN(new_n280_));
  XOR2_X1   g079(.A(G71gat), .B(G78gat), .Z(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n282_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT75), .Z(new_n284_));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285_));
  INV_X1    g084(.A(G1gat), .ZN(new_n286_));
  INV_X1    g085(.A(G8gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT14), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G1gat), .B(G8gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  NAND2_X1  g090(.A1(G231gat), .A2(G233gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n292_), .B(KEYINPUT74), .Z(new_n293_));
  XOR2_X1   g092(.A(new_n291_), .B(new_n293_), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n284_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT17), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G127gat), .B(G155gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G183gat), .B(G211gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n295_), .A2(new_n296_), .A3(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n302_), .B(KEYINPUT77), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n283_), .B(KEYINPUT69), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n294_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n301_), .B(KEYINPUT17), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n277_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT78), .ZN(new_n310_));
  XOR2_X1   g109(.A(G120gat), .B(G148gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G204gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT5), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT12), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n283_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n240_), .A2(new_n250_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT71), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n240_), .A2(new_n241_), .A3(new_n250_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n318_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n304_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n240_), .A2(new_n323_), .A3(new_n250_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n240_), .B2(new_n250_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(KEYINPUT12), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G230gat), .A2(G233gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n322_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n319_), .A2(new_n304_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(new_n330_), .B2(new_n324_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT70), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(KEYINPUT70), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n315_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT70), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n317_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n330_), .A2(new_n316_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n337_), .A2(new_n327_), .A3(new_n338_), .A4(new_n324_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n331_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n315_), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n341_), .A2(new_n333_), .A3(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n335_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT13), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n310_), .A2(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(KEYINPUT79), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT103), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT4), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G127gat), .B(G134gat), .ZN(new_n353_));
  INV_X1    g152(.A(G113gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G120gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT87), .Z(new_n359_));
  NAND2_X1  g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n360_), .B(KEYINPUT1), .Z(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT88), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT88), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n370_), .A3(new_n367_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n369_), .B(new_n371_), .C1(new_n367_), .C2(new_n365_), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n363_), .B(KEYINPUT3), .Z(new_n373_));
  OAI211_X1 g172(.A(new_n359_), .B(new_n360_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n366_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n357_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n366_), .A2(new_n374_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n356_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(KEYINPUT98), .A3(new_n378_), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n357_), .A2(new_n375_), .A3(KEYINPUT98), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n352_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n378_), .A2(KEYINPUT4), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n351_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G1gat), .B(G29gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G57gat), .B(G85gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  NAND3_X1  g187(.A1(new_n379_), .A2(new_n380_), .A3(new_n350_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n383_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n383_), .B2(new_n389_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT92), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G197gat), .B(G204gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT91), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n393_), .A2(KEYINPUT92), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(KEYINPUT92), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n395_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT21), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT21), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT23), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(G183gat), .B2(G190gat), .ZN(new_n408_));
  INV_X1    g207(.A(G169gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(new_n314_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT22), .B(G169gat), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(new_n314_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT25), .B(G183gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT96), .Z(new_n415_));
  XOR2_X1   g214(.A(KEYINPUT26), .B(G190gat), .Z(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n410_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n409_), .A2(new_n314_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT24), .A3(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n419_), .A2(KEYINPUT24), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n407_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n413_), .B1(new_n417_), .B2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n405_), .A2(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n424_), .A2(KEYINPUT97), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT20), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n424_), .B2(KEYINPUT97), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n428_), .B(KEYINPUT95), .Z(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT19), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n412_), .B(KEYINPUT84), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n408_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n416_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n434_), .A2(new_n414_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n435_), .A2(new_n422_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n405_), .A2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n425_), .A2(new_n427_), .A3(new_n431_), .A4(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n405_), .A2(new_n423_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n440_), .B(KEYINPUT20), .C1(new_n405_), .C2(new_n437_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n430_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT18), .B(G64gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(G92gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G8gat), .B(G36gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n444_), .B(new_n445_), .Z(new_n446_));
  AND3_X1   g245(.A1(new_n439_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT102), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT27), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n438_), .B1(new_n405_), .B2(new_n423_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n430_), .B1(new_n451_), .B2(new_n426_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n430_), .B2(new_n441_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n446_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n450_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n439_), .A2(new_n442_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT102), .B1(new_n456_), .B2(new_n454_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n449_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n446_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n450_), .B1(new_n447_), .B2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT94), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT93), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G22gat), .B(G50gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OR3_X1    g264(.A1(new_n377_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT89), .B1(new_n377_), .B2(KEYINPUT29), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n468_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n465_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n472_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(new_n464_), .A3(new_n470_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n463_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n377_), .A2(KEYINPUT29), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n402_), .A2(new_n404_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G228gat), .A2(G233gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(G228gat), .B(G233gat), .C1(new_n477_), .C2(new_n478_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G78gat), .B(G106gat), .Z(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n476_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n473_), .A2(new_n475_), .A3(new_n486_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n476_), .B2(new_n484_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n462_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n473_), .A2(new_n475_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n485_), .B1(new_n493_), .B2(new_n463_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n494_), .A2(KEYINPUT94), .A3(new_n490_), .A4(new_n488_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n433_), .A2(new_n496_), .A3(new_n436_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n498_), .A2(G71gat), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G71gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n437_), .A2(KEYINPUT30), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n497_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n357_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(G71gat), .B1(new_n498_), .B2(new_n499_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n501_), .A3(new_n497_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n356_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n509_));
  NAND2_X1  g308(.A1(G227gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G15gat), .B(G43gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(G99gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n511_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n508_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n504_), .A2(new_n507_), .A3(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n492_), .A2(new_n495_), .A3(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n516_), .A2(KEYINPUT86), .A3(new_n517_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT86), .B1(new_n516_), .B2(new_n517_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n392_), .B(new_n461_), .C1(new_n519_), .C2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n446_), .A2(KEYINPUT32), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n453_), .A2(new_n525_), .ZN(new_n526_));
  OAI221_X1 g325(.A(new_n526_), .B1(new_n456_), .B2(new_n525_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n447_), .A2(new_n459_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n379_), .A2(new_n380_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n351_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n381_), .A2(new_n382_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n388_), .B(new_n530_), .C1(new_n531_), .C2(new_n351_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n391_), .A2(KEYINPUT100), .A3(KEYINPUT33), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT100), .B1(new_n391_), .B2(KEYINPUT33), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n528_), .B(new_n532_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT101), .ZN(new_n536_));
  OR3_X1    g335(.A1(new_n391_), .A2(new_n536_), .A3(KEYINPUT33), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n536_), .B1(new_n391_), .B2(KEYINPUT33), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n527_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n492_), .A2(new_n495_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n522_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n524_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n291_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n205_), .A2(new_n209_), .A3(KEYINPUT80), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT80), .B1(new_n205_), .B2(new_n209_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT80), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n211_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n205_), .A2(new_n209_), .A3(KEYINPUT80), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n291_), .A3(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n548_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n213_), .A2(new_n545_), .A3(new_n210_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n554_), .B(KEYINPUT81), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT82), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT82), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n552_), .A2(new_n556_), .A3(new_n560_), .A4(new_n557_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(new_n409_), .ZN(new_n564_));
  INV_X1    g363(.A(G197gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(KEYINPUT83), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n562_), .B(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n349_), .B1(new_n544_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  AOI211_X1 g370(.A(KEYINPUT103), .B(new_n571_), .C1(new_n524_), .C2(new_n543_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n347_), .A2(KEYINPUT79), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n348_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n392_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n576_), .A2(KEYINPUT38), .A3(new_n286_), .A4(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n345_), .A2(new_n571_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n269_), .A2(new_n272_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n308_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n544_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G1gat), .B1(new_n585_), .B2(new_n392_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n348_), .A2(new_n286_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n587_), .B1(new_n588_), .B2(new_n392_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n578_), .A2(new_n586_), .A3(new_n589_), .ZN(G1324gat));
  INV_X1    g389(.A(new_n461_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n287_), .B1(new_n584_), .B2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT39), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n287_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n593_), .B1(new_n575_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT40), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(KEYINPUT40), .B(new_n593_), .C1(new_n575_), .C2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(G1325gat));
  INV_X1    g398(.A(G15gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n576_), .A2(new_n600_), .A3(new_n522_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n584_), .B2(new_n522_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT41), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(G1326gat));
  OAI21_X1  g403(.A(G22gat), .B1(new_n585_), .B2(new_n541_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT42), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n541_), .A2(G22gat), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n606_), .B1(new_n575_), .B2(new_n607_), .ZN(G1327gat));
  NOR2_X1   g407(.A1(new_n581_), .A2(new_n582_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n346_), .B(new_n609_), .C1(new_n570_), .C2(new_n572_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(G29gat), .B1(new_n611_), .B2(new_n577_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n544_), .A2(new_n613_), .A3(new_n277_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n544_), .B2(new_n277_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n579_), .B(new_n308_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT44), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n544_), .A2(new_n277_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT43), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n544_), .A2(new_n613_), .A3(new_n277_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n622_), .A2(KEYINPUT44), .A3(new_n579_), .A4(new_n308_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n392_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n612_), .B1(new_n625_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g425(.A(KEYINPUT46), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n461_), .A2(G36gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT45), .B1(new_n611_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT45), .ZN(new_n630_));
  NOR4_X1   g429(.A1(new_n610_), .A2(new_n630_), .A3(G36gat), .A4(new_n461_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n618_), .A2(new_n623_), .A3(new_n591_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G36gat), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n627_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n634_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT104), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(KEYINPUT46), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n642_), .ZN(G1329gat));
  INV_X1    g442(.A(KEYINPUT47), .ZN(new_n644_));
  INV_X1    g443(.A(new_n518_), .ZN(new_n645_));
  INV_X1    g444(.A(G43gat), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n618_), .A2(new_n623_), .A3(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n610_), .B2(new_n542_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT105), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n650_), .A2(KEYINPUT105), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n644_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(KEYINPUT47), .A3(new_n651_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1330gat));
  OAI21_X1  g456(.A(G50gat), .B1(new_n624_), .B2(new_n541_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n541_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n206_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT106), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n610_), .B2(new_n661_), .ZN(G1331gat));
  AOI21_X1  g461(.A(new_n569_), .B1(new_n524_), .B2(new_n543_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n663_), .A2(new_n345_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n664_));
  INV_X1    g463(.A(G57gat), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(new_n392_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n663_), .B(KEYINPUT107), .Z(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n346_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n310_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n668_), .A2(KEYINPUT108), .A3(new_n310_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n577_), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n666_), .B1(new_n673_), .B2(new_n665_), .ZN(G1332gat));
  OAI21_X1  g473(.A(G64gat), .B1(new_n664_), .B2(new_n461_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT48), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n672_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n461_), .A2(G64gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(G1333gat));
  OAI21_X1  g478(.A(G71gat), .B1(new_n664_), .B2(new_n542_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT49), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n522_), .A2(new_n501_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n677_), .B2(new_n682_), .ZN(G1334gat));
  OAI21_X1  g482(.A(G78gat), .B1(new_n664_), .B2(new_n541_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT50), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n541_), .A2(G78gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n677_), .B2(new_n686_), .ZN(G1335gat));
  NAND2_X1  g486(.A1(new_n622_), .A2(KEYINPUT109), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n345_), .A2(new_n571_), .A3(new_n308_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n620_), .A2(new_n691_), .A3(new_n621_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n688_), .A2(new_n690_), .A3(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(G85gat), .A3(new_n577_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n668_), .A2(new_n609_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(new_n392_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n696_), .B2(G85gat), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(G1336gat));
  NAND3_X1  g497(.A1(new_n693_), .A2(G92gat), .A3(new_n591_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n695_), .A2(new_n461_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G92gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(G1337gat));
  NOR2_X1   g501(.A1(new_n645_), .A2(new_n247_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n668_), .A2(new_n609_), .A3(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n688_), .A2(new_n522_), .A3(new_n690_), .A4(new_n692_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(KEYINPUT110), .A3(G99gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT110), .B1(new_n705_), .B2(G99gat), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT111), .B(new_n704_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT51), .ZN(new_n710_));
  INV_X1    g509(.A(new_n708_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n706_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n712_), .A2(KEYINPUT111), .A3(new_n713_), .A4(new_n704_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(new_n714_), .ZN(G1338gat));
  NAND3_X1  g514(.A1(new_n622_), .A2(new_n659_), .A3(new_n690_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT52), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(G106gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G106gat), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n541_), .A2(G106gat), .ZN(new_n720_));
  OAI22_X1  g519(.A1(new_n718_), .A2(new_n719_), .B1(new_n695_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT53), .ZN(G1339gat));
  XOR2_X1   g521(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT113), .Z(new_n724_));
  NOR3_X1   g523(.A1(new_n277_), .A2(new_n569_), .A3(new_n308_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n346_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n723_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(KEYINPUT113), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n725_), .A2(new_n346_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n332_), .A2(new_n334_), .A3(new_n315_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n569_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n733_), .B1(new_n322_), .B2(new_n326_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n240_), .A2(new_n323_), .A3(new_n250_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n330_), .B2(new_n316_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(KEYINPUT114), .A3(new_n337_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n737_), .A3(new_n328_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n322_), .A2(new_n326_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n739_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n327_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n736_), .A2(new_n337_), .A3(KEYINPUT55), .A4(new_n327_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n339_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n738_), .A2(new_n740_), .A3(new_n743_), .A4(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n342_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(KEYINPUT56), .A3(new_n342_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n732_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n555_), .A2(new_n567_), .A3(new_n559_), .A4(new_n561_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n557_), .ZN(new_n753_));
  OAI211_X1 g552(.A(KEYINPUT116), .B(new_n566_), .C1(new_n553_), .C2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n753_), .B1(new_n548_), .B2(new_n552_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n567_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n552_), .A2(new_n556_), .A3(new_n753_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n752_), .A2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT117), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n344_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n581_), .B1(new_n751_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT56), .B1(new_n746_), .B2(new_n342_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n746_), .A2(KEYINPUT56), .A3(new_n342_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n343_), .A2(new_n768_), .A3(new_n761_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n760_), .B(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT118), .B1(new_n731_), .B2(new_n771_), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n766_), .A2(new_n767_), .B1(new_n769_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n768_), .B1(new_n343_), .B2(new_n761_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n731_), .A2(new_n771_), .A3(KEYINPUT118), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(KEYINPUT58), .C1(new_n766_), .C2(new_n767_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n277_), .A3(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT57), .B(new_n581_), .C1(new_n751_), .C2(new_n762_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n765_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n308_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n730_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n591_), .A2(new_n392_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n519_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G113gat), .B1(new_n788_), .B2(new_n569_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n783_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n782_), .A2(KEYINPUT120), .A3(new_n308_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n730_), .A3(new_n792_), .ZN(new_n793_));
  XOR2_X1   g592(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n786_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n787_), .A2(KEYINPUT59), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n354_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n789_), .B1(new_n798_), .B2(new_n569_), .ZN(G1340gat));
  OAI21_X1  g598(.A(G120gat), .B1(new_n797_), .B2(new_n346_), .ZN(new_n800_));
  INV_X1    g599(.A(G120gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n346_), .B2(KEYINPUT60), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n801_), .A2(KEYINPUT60), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n784_), .A2(new_n786_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT121), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n800_), .A2(new_n805_), .ZN(G1341gat));
  AOI21_X1  g605(.A(G127gat), .B1(new_n788_), .B2(new_n582_), .ZN(new_n807_));
  OAI21_X1  g606(.A(G127gat), .B1(new_n308_), .B2(KEYINPUT122), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n795_), .A2(new_n796_), .A3(new_n808_), .ZN(new_n809_));
  OR2_X1    g608(.A1(KEYINPUT122), .A2(G127gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n807_), .B1(new_n809_), .B2(new_n810_), .ZN(G1342gat));
  INV_X1    g610(.A(new_n581_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G134gat), .B1(new_n788_), .B2(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n795_), .A2(new_n277_), .A3(new_n796_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g614(.A1(new_n784_), .A2(new_n523_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n785_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n816_), .A2(new_n571_), .A3(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT123), .B(G141gat), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1344gat));
  INV_X1    g619(.A(new_n816_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(new_n345_), .A3(new_n785_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(G148gat), .ZN(G1345gat));
  NOR3_X1   g622(.A1(new_n816_), .A2(new_n308_), .A3(new_n817_), .ZN(new_n824_));
  XOR2_X1   g623(.A(KEYINPUT61), .B(G155gat), .Z(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(G1346gat));
  NOR3_X1   g625(.A1(new_n816_), .A2(new_n581_), .A3(new_n817_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n821_), .A2(new_n277_), .A3(new_n785_), .ZN(new_n828_));
  MUX2_X1   g627(.A(new_n827_), .B(new_n828_), .S(G162gat), .Z(G1347gat));
  NOR2_X1   g628(.A1(new_n461_), .A2(new_n577_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n522_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n659_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n793_), .A2(new_n569_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G169gat), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n837_));
  INV_X1    g636(.A(new_n411_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n836_), .B(new_n837_), .C1(new_n838_), .C2(new_n833_), .ZN(G1348gat));
  NAND3_X1  g638(.A1(new_n793_), .A2(new_n345_), .A3(new_n832_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n314_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n659_), .B1(new_n730_), .B2(new_n783_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n346_), .A2(new_n314_), .A3(new_n831_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n841_), .A2(KEYINPUT124), .A3(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1349gat));
  NOR2_X1   g648(.A1(new_n831_), .A2(new_n308_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G183gat), .B1(new_n842_), .B2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n793_), .A2(new_n832_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n582_), .A2(new_n415_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1350gat));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n277_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G190gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n852_), .A2(new_n812_), .A3(new_n434_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1351gat));
  NAND3_X1  g657(.A1(new_n784_), .A2(new_n523_), .A3(new_n830_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n571_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(KEYINPUT125), .A3(new_n565_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT125), .B(G197gat), .Z(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n860_), .B2(new_n862_), .ZN(G1352gat));
  AND3_X1   g662(.A1(new_n784_), .A2(new_n523_), .A3(new_n830_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n345_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g665(.A(KEYINPUT126), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n308_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n864_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n868_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT126), .B1(new_n859_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n873_));
  INV_X1    g672(.A(G211gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n869_), .A2(new_n871_), .A3(new_n873_), .A4(new_n874_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1354gat));
  AOI21_X1  g677(.A(G218gat), .B1(new_n864_), .B2(new_n812_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n277_), .A2(G218gat), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n880_), .B(KEYINPUT127), .Z(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n864_), .B2(new_n881_), .ZN(G1355gat));
endmodule


