//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n922_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT82), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n203_), .B1(G169gat), .B2(G176gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT96), .B(KEYINPUT24), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT23), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n202_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n206_), .B(new_n212_), .C1(new_n213_), .C2(new_n205_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT22), .B(G169gat), .Z(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT97), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n215_), .B(new_n216_), .C1(new_n218_), .C2(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G204gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT91), .B1(new_n221_), .B2(G197gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(G197gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n221_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT21), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G211gat), .B(G218gat), .Z(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n223_), .B(KEYINPUT92), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n229_), .B1(G197gat), .B2(new_n221_), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n226_), .B(new_n228_), .C1(new_n230_), .C2(KEYINPUT21), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT21), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(new_n227_), .B2(KEYINPUT93), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n230_), .B(new_n233_), .C1(KEYINPUT93), .C2(new_n227_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n220_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT83), .B1(KEYINPUT84), .B2(G169gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT22), .ZN(new_n238_));
  INV_X1    g037(.A(G176gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT22), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(KEYINPUT84), .A3(G169gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT83), .B1(new_n240_), .B2(G169gat), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n238_), .A2(new_n239_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n215_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT85), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n216_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n204_), .A2(KEYINPUT24), .ZN(new_n247_));
  INV_X1    g046(.A(new_n203_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n247_), .B(new_n212_), .C1(KEYINPUT24), .C2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n236_), .B(KEYINPUT20), .C1(new_n250_), .C2(new_n235_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT19), .Z(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT95), .Z(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT20), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n250_), .B2(new_n235_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n257_), .B(new_n253_), .C1(new_n235_), .C2(new_n220_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G8gat), .B(G36gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT18), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(G64gat), .ZN(new_n262_));
  INV_X1    g061(.A(G92gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n259_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n255_), .A2(new_n258_), .A3(new_n264_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT27), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n251_), .A2(new_n254_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT103), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n220_), .A2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n231_), .A2(new_n234_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n214_), .A2(KEYINPUT103), .A3(new_n219_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n253_), .B1(new_n276_), .B2(new_n257_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n265_), .B1(new_n271_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(KEYINPUT27), .A3(new_n267_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n270_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G141gat), .A2(G148gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G141gat), .A2(G148gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT1), .Z(new_n284_));
  NOR2_X1   g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT89), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n282_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n286_), .A2(new_n283_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n281_), .B(KEYINPUT2), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n282_), .B1(KEYINPUT90), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT90), .B(KEYINPUT3), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n289_), .B(new_n291_), .C1(new_n282_), .C2(new_n292_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n281_), .A2(new_n287_), .B1(new_n288_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(KEYINPUT28), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(KEYINPUT28), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n298_), .A2(G228gat), .A3(G233gat), .A4(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  INV_X1    g100(.A(G228gat), .ZN(new_n302_));
  INV_X1    g101(.A(G233gat), .ZN(new_n303_));
  OAI22_X1  g102(.A1(new_n301_), .A2(new_n297_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G22gat), .B(G50gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n300_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n294_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n274_), .B1(new_n309_), .B2(KEYINPUT29), .ZN(new_n310_));
  XOR2_X1   g109(.A(G78gat), .B(G106gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT94), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n310_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n306_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n308_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n313_), .B1(new_n317_), .B2(new_n307_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT105), .B1(new_n280_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G127gat), .B(G134gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT86), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G113gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n321_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G113gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G120gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n323_), .A2(new_n327_), .A3(G120gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT31), .Z(new_n333_));
  INV_X1    g132(.A(G43gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n250_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G71gat), .B(G99gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT30), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G227gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G15gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n337_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n335_), .B(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n333_), .B1(new_n341_), .B2(KEYINPUT87), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(KEYINPUT87), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n294_), .A2(KEYINPUT98), .ZN(new_n345_));
  INV_X1    g144(.A(new_n331_), .ZN(new_n346_));
  AOI21_X1  g145(.A(G120gat), .B1(new_n323_), .B2(new_n327_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n330_), .A2(KEYINPUT98), .A3(new_n294_), .A4(new_n331_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(KEYINPUT4), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n332_), .A2(new_n351_), .A3(new_n309_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G57gat), .B(G85gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NOR2_X1   g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n354_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n366_), .B2(new_n357_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n316_), .A2(new_n318_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT105), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n370_), .A2(new_n270_), .A3(new_n371_), .A4(new_n279_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n320_), .A2(new_n344_), .A3(new_n369_), .A4(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT106), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT100), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n376_), .B1(new_n367_), .B2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n359_), .A2(KEYINPUT100), .A3(KEYINPUT33), .A4(new_n364_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n364_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n348_), .A2(new_n349_), .A3(new_n355_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n381_), .B(new_n382_), .C1(new_n353_), .C2(new_n355_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n266_), .A2(new_n267_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n367_), .A2(KEYINPUT101), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT101), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n386_), .B(new_n364_), .C1(new_n366_), .C2(new_n357_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n377_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n380_), .A2(new_n384_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT102), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n271_), .B2(new_n277_), .ZN(new_n392_));
  OAI221_X1 g191(.A(new_n392_), .B1(new_n259_), .B2(new_n391_), .C1(new_n365_), .C2(new_n368_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT102), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n380_), .A2(new_n384_), .A3(new_n388_), .A4(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n370_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT104), .ZN(new_n398_));
  INV_X1    g197(.A(new_n280_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n369_), .A3(new_n319_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT104), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n396_), .A2(new_n401_), .A3(new_n370_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n344_), .B(KEYINPUT88), .Z(new_n404_));
  AOI21_X1  g203(.A(new_n375_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G99gat), .ZN(new_n406_));
  INV_X1    g205(.A(G106gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT65), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT7), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n408_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n406_), .B(new_n407_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT64), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT64), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT6), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G99gat), .A2(G106gat), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n416_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n413_), .B(new_n414_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G85gat), .B(G92gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT67), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G85gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n263_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G85gat), .A2(G92gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(KEYINPUT67), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n422_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT8), .B1(new_n430_), .B2(KEYINPUT66), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n422_), .B(new_n430_), .C1(KEYINPUT66), .C2(KEYINPUT8), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n420_), .A2(new_n421_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT10), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n436_), .A2(G99gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n406_), .A2(KEYINPUT10), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n407_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n427_), .A2(KEYINPUT9), .A3(new_n428_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n428_), .A2(KEYINPUT9), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n433_), .A2(new_n434_), .A3(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(G57gat), .A2(G64gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(G57gat), .A2(G64gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT11), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n452_));
  INV_X1    g251(.A(G71gat), .ZN(new_n453_));
  INV_X1    g252(.A(G78gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n454_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n452_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G57gat), .ZN(new_n459_));
  INV_X1    g258(.A(G64gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G57gat), .A2(G64gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n449_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n455_), .ZN(new_n464_));
  AND4_X1   g263(.A1(new_n452_), .A2(new_n463_), .A3(new_n457_), .A4(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n451_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(new_n452_), .A3(new_n457_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n464_), .A3(new_n457_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT68), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n469_), .A3(new_n450_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT12), .B1(new_n445_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n445_), .A2(new_n471_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT12), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n466_), .B2(new_n470_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n435_), .A2(new_n441_), .A3(KEYINPUT69), .A4(new_n443_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT69), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n440_), .B(new_n439_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n442_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n433_), .A2(new_n434_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n476_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT70), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G230gat), .A2(G233gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n477_), .A2(new_n480_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(new_n434_), .A3(new_n433_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(KEYINPUT70), .A3(new_n476_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n474_), .A2(new_n485_), .A3(new_n486_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n473_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n445_), .A2(new_n471_), .ZN(new_n492_));
  OAI211_X1 g291(.A(G230gat), .B(G233gat), .C1(new_n491_), .C2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G120gat), .B(G148gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT5), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G176gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G204gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n490_), .A2(new_n493_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n501_), .A2(KEYINPUT13), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(KEYINPUT13), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  INV_X1    g304(.A(G50gat), .ZN(new_n506_));
  INV_X1    g305(.A(G29gat), .ZN(new_n507_));
  INV_X1    g306(.A(G36gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT72), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT72), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n513_), .A3(new_n510_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n334_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n334_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n506_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n512_), .A2(new_n514_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(G43gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(G50gat), .A3(new_n515_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G8gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT79), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G15gat), .ZN(new_n527_));
  INV_X1    g326(.A(G22gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G15gat), .A2(G22gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G1gat), .A2(G8gat), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n529_), .A2(new_n530_), .B1(KEYINPUT14), .B2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n526_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n523_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n522_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n505_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT81), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n518_), .A2(new_n521_), .A3(KEYINPUT15), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT15), .B1(new_n518_), .B2(new_n521_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n505_), .B(new_n534_), .C1(new_n541_), .C2(new_n533_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n534_), .A2(new_n536_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n505_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n538_), .B1(new_n546_), .B2(KEYINPUT81), .ZN(new_n547_));
  XOR2_X1   g346(.A(G113gat), .B(G141gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(G169gat), .ZN(new_n549_));
  INV_X1    g348(.A(G197gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT81), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n545_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n535_), .A2(new_n522_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT15), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n522_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n518_), .A2(new_n521_), .A3(KEYINPUT15), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n556_), .B1(new_n560_), .B2(new_n535_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n537_), .B1(new_n561_), .B2(new_n505_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n555_), .B(new_n552_), .C1(new_n562_), .C2(new_n554_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n553_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n504_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n405_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n488_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT73), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n560_), .A2(KEYINPUT73), .A3(new_n488_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT34), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(KEYINPUT35), .ZN(new_n575_));
  INV_X1    g374(.A(new_n445_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(new_n523_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n571_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(KEYINPUT35), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT71), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT75), .ZN(new_n583_));
  INV_X1    g382(.A(new_n569_), .ZN(new_n584_));
  OAI221_X1 g383(.A(new_n580_), .B1(KEYINPUT35), .B2(new_n574_), .C1(new_n445_), .C2(new_n522_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n583_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n577_), .A2(new_n569_), .A3(KEYINPUT75), .A4(new_n580_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT74), .ZN(new_n591_));
  INV_X1    g390(.A(G134gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(G162gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT36), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n589_), .A2(new_n595_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n581_), .A2(new_n578_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT76), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  AND4_X1   g398(.A1(KEYINPUT76), .A2(new_n582_), .A3(new_n588_), .A4(new_n598_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n596_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT37), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT76), .ZN(new_n603_));
  INV_X1    g402(.A(new_n598_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n603_), .B1(new_n589_), .B2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n597_), .A2(KEYINPUT76), .A3(new_n598_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT77), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n589_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n597_), .A2(KEYINPUT77), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n595_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n607_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT78), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n602_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n602_), .B2(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n533_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n471_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT17), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT16), .ZN(new_n622_));
  INV_X1    g421(.A(G183gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(G211gat), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n619_), .A2(new_n620_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT80), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n625_), .B(KEYINPUT17), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n619_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n615_), .A2(new_n616_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n568_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT107), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n633_), .A2(G1gat), .A3(new_n369_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT38), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n607_), .A2(new_n611_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n630_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n568_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n369_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n634_), .A2(KEYINPUT38), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n641_), .A3(new_n642_), .ZN(G1324gat));
  NAND2_X1  g442(.A1(new_n403_), .A2(new_n404_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n375_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n646_), .A2(new_n566_), .A3(new_n280_), .A4(new_n638_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT108), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n568_), .A2(KEYINPUT108), .A3(new_n280_), .A4(new_n638_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(G8gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n649_), .A2(new_n650_), .A3(new_n653_), .A4(G8gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n399_), .A2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n633_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n655_), .B(KEYINPUT40), .C1(new_n633_), .C2(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1325gat));
  INV_X1    g460(.A(new_n404_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n527_), .B1(new_n639_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  INV_X1    g463(.A(new_n633_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n527_), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1326gat));
  XNOR2_X1  g466(.A(new_n319_), .B(KEYINPUT109), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n528_), .B1(new_n639_), .B2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT42), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n665_), .A2(new_n528_), .A3(new_n669_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(new_n630_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n636_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n568_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n369_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n507_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n615_), .A2(new_n616_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n646_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n405_), .B2(new_n680_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n566_), .A3(new_n630_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n684_), .A2(KEYINPUT44), .A3(new_n566_), .A4(new_n630_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n677_), .A3(new_n688_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n689_), .A2(KEYINPUT110), .A3(G29gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT110), .B1(new_n689_), .B2(G29gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n678_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  AOI211_X1 g492(.A(new_n567_), .B(new_n674_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n399_), .B1(new_n694_), .B2(KEYINPUT44), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n508_), .B1(new_n695_), .B2(new_n687_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n676_), .A2(new_n508_), .A3(new_n280_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n693_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n687_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n688_), .A2(new_n280_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G36gat), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n697_), .B(KEYINPUT45), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(KEYINPUT46), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n705_), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n687_), .A2(G43gat), .A3(new_n344_), .A4(new_n688_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n676_), .A2(new_n662_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n334_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT47), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1330gat));
  NAND2_X1  g513(.A1(new_n688_), .A2(new_n319_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G50gat), .B1(new_n701_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n669_), .A2(new_n506_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT111), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n676_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(new_n504_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n565_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n405_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(new_n631_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n677_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n725_), .A2(new_n638_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n369_), .A2(new_n459_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(G1332gat));
  AOI21_X1  g529(.A(new_n460_), .B1(new_n728_), .B2(new_n280_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT48), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n726_), .A2(new_n460_), .A3(new_n280_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1333gat));
  AOI21_X1  g533(.A(new_n453_), .B1(new_n728_), .B2(new_n662_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT49), .Z(new_n736_));
  NAND3_X1  g535(.A1(new_n726_), .A2(new_n453_), .A3(new_n662_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1334gat));
  AOI21_X1  g537(.A(new_n454_), .B1(new_n728_), .B2(new_n669_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT50), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n726_), .A2(new_n454_), .A3(new_n669_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1335gat));
  AND2_X1   g541(.A1(new_n725_), .A2(new_n675_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n677_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n724_), .A2(new_n674_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT112), .B1(new_n684_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747_));
  INV_X1    g546(.A(new_n745_), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n747_), .B(new_n748_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n746_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n369_), .A2(new_n426_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n744_), .B1(new_n750_), .B2(new_n751_), .ZN(G1336gat));
  AOI21_X1  g551(.A(G92gat), .B1(new_n743_), .B2(new_n280_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n399_), .A2(new_n263_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n750_), .B2(new_n754_), .ZN(G1337gat));
  OAI211_X1 g554(.A(new_n743_), .B(new_n344_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n746_), .A2(new_n749_), .A3(new_n404_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n406_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT51), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n756_), .C1(new_n757_), .C2(new_n406_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1338gat));
  NAND3_X1  g561(.A1(new_n684_), .A2(new_n319_), .A3(new_n745_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G106gat), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(KEYINPUT113), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n743_), .A2(new_n407_), .A3(new_n319_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n765_), .A2(KEYINPUT113), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(KEYINPUT113), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n763_), .A2(G106gat), .A3(new_n768_), .A4(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n766_), .A2(new_n767_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n766_), .A2(new_n773_), .A3(new_n767_), .A4(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  NAND2_X1  g574(.A1(new_n561_), .A2(new_n544_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n543_), .A2(new_n505_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n551_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT116), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n776_), .A2(new_n777_), .A3(new_n780_), .A4(new_n551_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n563_), .A2(new_n779_), .A3(new_n498_), .A4(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n474_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(G230gat), .A3(G233gat), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n488_), .A2(KEYINPUT70), .A3(new_n476_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT70), .B1(new_n488_), .B2(new_n476_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n790_), .A2(KEYINPUT55), .A3(new_n486_), .A4(new_n474_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n490_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n490_), .B2(new_n794_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n792_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n785_), .B1(new_n797_), .B2(new_n497_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n490_), .A2(new_n794_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT115), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n490_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n800_), .A2(new_n787_), .A3(new_n791_), .A4(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n497_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n798_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n784_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n784_), .A2(new_n805_), .A3(KEYINPUT58), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n808_), .B(new_n809_), .C1(new_n616_), .C2(new_n615_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n498_), .B1(new_n553_), .B2(new_n564_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n803_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n803_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n563_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(new_n501_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n637_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n819_), .A2(KEYINPUT117), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n811_), .B1(new_n798_), .B2(new_n804_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n636_), .B1(new_n822_), .B2(new_n817_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT57), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n810_), .B1(new_n821_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT119), .B(new_n810_), .C1(new_n821_), .C2(new_n825_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n630_), .A3(new_n829_), .ZN(new_n830_));
  NOR4_X1   g629(.A1(new_n615_), .A2(new_n616_), .A3(new_n722_), .A4(new_n630_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n721_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT54), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n631_), .A2(new_n834_), .A3(new_n565_), .A4(new_n721_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT114), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n831_), .A2(new_n837_), .A3(new_n834_), .A4(new_n721_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n830_), .A2(new_n839_), .ZN(new_n840_));
  AND4_X1   g639(.A1(new_n677_), .A2(new_n320_), .A3(new_n344_), .A4(new_n372_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842_), .B2(new_n722_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n826_), .A2(new_n630_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n839_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n844_), .A3(new_n841_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n565_), .A2(new_n326_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n843_), .B1(new_n850_), .B2(new_n851_), .ZN(G1340gat));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n721_), .B2(G120gat), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n842_), .B(new_n854_), .C1(new_n853_), .C2(G120gat), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(G120gat), .B1(new_n849_), .B2(new_n721_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1341gat));
  AOI21_X1  g658(.A(G127gat), .B1(new_n842_), .B2(new_n674_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n674_), .A2(G127gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n850_), .B2(new_n861_), .ZN(G1342gat));
  AOI21_X1  g661(.A(G134gat), .B1(new_n842_), .B2(new_n637_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n680_), .A2(new_n592_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n850_), .B2(new_n864_), .ZN(G1343gat));
  AOI21_X1  g664(.A(new_n662_), .B1(new_n830_), .B2(new_n839_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n866_), .A2(new_n677_), .A3(new_n399_), .A4(new_n319_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n565_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n721_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT121), .B(G148gat), .Z(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n867_), .A2(new_n630_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT122), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n873_), .B(new_n875_), .ZN(G1346gat));
  OR3_X1    g675(.A1(new_n867_), .A2(G162gat), .A3(new_n636_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878_));
  OAI21_X1  g677(.A(G162gat), .B1(new_n867_), .B2(new_n680_), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n399_), .A2(new_n677_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n662_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n847_), .A2(new_n668_), .A3(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G169gat), .B1(new_n886_), .B2(new_n565_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n565_), .A2(new_n218_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT124), .ZN(new_n891_));
  OAI22_X1  g690(.A1(new_n888_), .A2(new_n889_), .B1(new_n886_), .B2(new_n891_), .ZN(G1348gat));
  NAND2_X1  g691(.A1(new_n840_), .A2(new_n370_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n840_), .A2(KEYINPUT125), .A3(new_n370_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n895_), .A2(G176gat), .A3(new_n885_), .A4(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT126), .B1(new_n897_), .B2(new_n721_), .ZN(new_n898_));
  AOI21_X1  g697(.A(KEYINPUT125), .B1(new_n840_), .B2(new_n370_), .ZN(new_n899_));
  AOI211_X1 g698(.A(new_n894_), .B(new_n319_), .C1(new_n830_), .C2(new_n839_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n884_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(G176gat), .A4(new_n504_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n239_), .B1(new_n886_), .B2(new_n721_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n898_), .A2(new_n903_), .A3(new_n904_), .ZN(G1349gat));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  AOI21_X1  g705(.A(G183gat), .B1(new_n901_), .B2(new_n674_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n886_), .A2(new_n207_), .A3(new_n630_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n895_), .A2(new_n885_), .A3(new_n896_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n623_), .B1(new_n910_), .B2(new_n630_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n908_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(KEYINPUT127), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n909_), .A2(new_n913_), .ZN(G1350gat));
  INV_X1    g713(.A(new_n886_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n208_), .A3(new_n637_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G190gat), .B1(new_n886_), .B2(new_n680_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1351gat));
  AND3_X1   g717(.A1(new_n866_), .A2(new_n319_), .A3(new_n883_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n722_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n504_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g722(.A1(new_n919_), .A2(new_n674_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n924_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT63), .B(G211gat), .Z(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n924_), .B2(new_n926_), .ZN(G1354gat));
  AOI21_X1  g726(.A(G218gat), .B1(new_n919_), .B2(new_n637_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n681_), .A2(G218gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n919_), .B2(new_n929_), .ZN(G1355gat));
endmodule


