//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT13), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT7), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(new_n207_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n205_), .A2(new_n208_), .A3(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G85gat), .B(G92gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT8), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(new_n210_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT65), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n207_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n205_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n214_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n216_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT9), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n229_), .B(new_n232_), .C1(new_n214_), .C2(new_n231_), .ZN(new_n233_));
  OR2_X1    g032(.A1(G85gat), .A2(G92gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n231_), .B1(new_n234_), .B2(new_n230_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n232_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT64), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n217_), .A2(new_n210_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n220_), .A2(new_n222_), .A3(new_n207_), .ZN(new_n240_));
  INV_X1    g039(.A(G99gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT10), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT10), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G99gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(G106gat), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n239_), .A2(new_n240_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n238_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n238_), .B2(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n228_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G57gat), .B(G64gat), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT11), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(KEYINPUT11), .ZN(new_n253_));
  XOR2_X1   g052(.A(G71gat), .B(G78gat), .Z(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n253_), .A2(new_n254_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(KEYINPUT12), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n238_), .A2(new_n246_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n228_), .A2(new_n261_), .A3(new_n257_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n215_), .A2(KEYINPUT8), .B1(new_n224_), .B2(new_n226_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n238_), .A2(new_n246_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n258_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n259_), .A2(new_n260_), .A3(new_n262_), .A4(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n262_), .A2(new_n265_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(G230gat), .A3(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(G204gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT5), .ZN(new_n274_));
  INV_X1    g073(.A(G176gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n268_), .A2(new_n270_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n268_), .A2(new_n270_), .A3(KEYINPUT69), .A4(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n268_), .A2(new_n270_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT68), .ZN(new_n283_));
  INV_X1    g082(.A(new_n276_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n268_), .A2(new_n285_), .A3(new_n270_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n281_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n281_), .B2(new_n287_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n203_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n281_), .A2(new_n287_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT70), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n281_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT13), .A3(new_n294_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n291_), .A2(new_n295_), .A3(KEYINPUT71), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT71), .B1(new_n291_), .B2(new_n295_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G29gat), .B(G36gat), .ZN(new_n299_));
  INV_X1    g098(.A(G43gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G50gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT15), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G15gat), .B(G22gat), .ZN(new_n305_));
  INV_X1    g104(.A(G8gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G8gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G229gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n301_), .B(G50gat), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n311_), .B(new_n312_), .C1(new_n313_), .C2(new_n310_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n310_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(G229gat), .A3(G233gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G113gat), .B(G141gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(G169gat), .B(G197gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n314_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G226gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT19), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT20), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT92), .ZN(new_n331_));
  XOR2_X1   g130(.A(G211gat), .B(G218gat), .Z(new_n332_));
  INV_X1    g131(.A(G197gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT88), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT88), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G197gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT89), .B1(new_n333_), .B2(G204gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT89), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(new_n272_), .A3(G197gat), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n337_), .A2(G204gat), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n332_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n340_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT88), .B(G197gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n344_), .B(new_n342_), .C1(new_n272_), .C2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT21), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n331_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n332_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n344_), .B1(new_n272_), .B2(new_n345_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(KEYINPUT91), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n353_), .A3(KEYINPUT92), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n332_), .B1(new_n341_), .B2(new_n352_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT90), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G197gat), .A2(G204gat), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT21), .B(new_n357_), .C1(new_n345_), .C2(G204gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n344_), .B(new_n352_), .C1(new_n272_), .C2(new_n345_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n349_), .A3(new_n358_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT90), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n348_), .A2(new_n354_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G169gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n275_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT23), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(G183gat), .A3(G190gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G183gat), .ZN(new_n374_));
  INV_X1    g173(.A(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n368_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT25), .B(G183gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT26), .B(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT82), .ZN(new_n382_));
  INV_X1    g181(.A(G169gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n275_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(KEYINPUT24), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(KEYINPUT24), .A3(new_n366_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n379_), .A2(new_n380_), .A3(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n382_), .A2(new_n386_), .A3(new_n387_), .A4(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n378_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n330_), .B1(new_n363_), .B2(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n343_), .A2(new_n347_), .A3(new_n331_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT92), .B1(new_n351_), .B2(new_n353_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n356_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n361_), .A2(KEYINPUT90), .ZN(new_n397_));
  OAI22_X1  g196(.A1(new_n394_), .A2(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(KEYINPUT95), .A2(KEYINPUT24), .ZN(new_n399_));
  NAND2_X1  g198(.A1(KEYINPUT95), .A2(KEYINPUT24), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n384_), .A3(new_n366_), .A4(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT96), .B1(new_n381_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n384_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n381_), .A2(KEYINPUT96), .A3(new_n401_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n377_), .A2(KEYINPUT97), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT97), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n373_), .A2(new_n409_), .A3(new_n376_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n368_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n398_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n329_), .B1(new_n393_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n330_), .B1(new_n398_), .B2(new_n391_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n348_), .A2(new_n354_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n359_), .A2(new_n362_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n367_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n381_), .A2(KEYINPUT96), .A3(new_n401_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(new_n402_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n422_), .B2(new_n405_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n418_), .A2(new_n419_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT98), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT98), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n363_), .A2(new_n426_), .A3(new_n423_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n417_), .A2(new_n425_), .A3(new_n329_), .A4(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT99), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n428_), .A2(new_n429_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n416_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT18), .B(G64gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G92gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n424_), .A2(KEYINPUT98), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT20), .B1(new_n363_), .B2(new_n392_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n441_), .A2(KEYINPUT99), .A3(new_n329_), .A4(new_n425_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n428_), .A2(new_n429_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(new_n416_), .A3(new_n436_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT0), .B(G57gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G85gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(G1gat), .B(G29gat), .Z(new_n448_));
  XOR2_X1   g247(.A(new_n447_), .B(new_n448_), .Z(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G113gat), .ZN(new_n451_));
  INV_X1    g250(.A(G127gat), .ZN(new_n452_));
  INV_X1    g251(.A(G134gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G127gat), .A2(G134gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n451_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(new_n451_), .A3(new_n455_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n457_), .A2(G120gat), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(G120gat), .B1(new_n457_), .B2(new_n458_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462_));
  OR2_X1    g261(.A1(G155gat), .A2(G162gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(G155gat), .A2(G162gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G155gat), .A2(G162gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT86), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  NOR4_X1   g269(.A1(KEYINPUT85), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT3), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G141gat), .A2(G148gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n470_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(new_n473_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n465_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT84), .B1(new_n465_), .B2(KEYINPUT1), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT1), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n468_), .B1(new_n467_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n483_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n462_), .B1(new_n480_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n473_), .A2(new_n474_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT3), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n473_), .A2(new_n474_), .A3(new_n472_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n479_), .A3(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(new_n469_), .A3(new_n466_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n485_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n465_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n488_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n482_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(KEYINPUT87), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n461_), .B1(new_n490_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n499_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n502_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G225gat), .A2(G233gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n450_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n459_), .A2(new_n460_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n480_), .A2(new_n489_), .A3(new_n462_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT87), .B1(new_n495_), .B2(new_n499_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n502_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n461_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(KEYINPUT4), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n515_), .B(new_n508_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n505_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n507_), .A2(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n501_), .A2(new_n503_), .A3(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n506_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT100), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT100), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n514_), .A2(new_n522_), .A3(new_n506_), .A4(new_n516_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n504_), .A2(new_n505_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n521_), .A2(new_n523_), .A3(new_n450_), .A4(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT33), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n438_), .A2(new_n445_), .A3(new_n518_), .A4(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n521_), .A2(new_n524_), .A3(new_n523_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n449_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n525_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n418_), .A2(new_n392_), .A3(new_n419_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n414_), .A2(KEYINPUT20), .A3(new_n329_), .A4(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT102), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT101), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n423_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n413_), .A2(KEYINPUT101), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n535_), .A2(new_n363_), .A3(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n328_), .B1(new_n537_), .B2(new_n440_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT102), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n393_), .A2(new_n539_), .A3(new_n414_), .A4(new_n329_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n533_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n436_), .A2(KEYINPUT32), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n530_), .A2(new_n544_), .ZN(new_n545_));
  AOI211_X1 g344(.A(new_n415_), .B(new_n543_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT103), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n444_), .A2(new_n416_), .A3(new_n542_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT103), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n530_), .A4(new_n544_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n527_), .A2(new_n547_), .A3(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G15gat), .B(G43gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT31), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n391_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G71gat), .B(G99gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n508_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G227gat), .A2(G233gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT30), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n461_), .B(new_n556_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(new_n559_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n555_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n559_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n554_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n564_), .A2(KEYINPUT83), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT83), .B1(new_n564_), .B2(new_n567_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT29), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n490_), .A2(new_n572_), .A3(new_n500_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G22gat), .B(G50gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT28), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT93), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n576_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G78gat), .B(G106gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n581_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n577_), .A2(new_n579_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n490_), .A2(new_n500_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n585_), .A2(KEYINPUT29), .B1(G228gat), .B2(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n398_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n512_), .A2(new_n572_), .ZN(new_n588_));
  OAI211_X1 g387(.A(G228gat), .B(G233gat), .C1(new_n363_), .C2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT94), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n582_), .B(new_n584_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n582_), .A2(new_n584_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n593_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(new_n591_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n571_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n551_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n438_), .A2(new_n445_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT27), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n570_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n564_), .A2(new_n567_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n594_), .A2(new_n597_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n530_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n541_), .A2(new_n437_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n445_), .A2(KEYINPUT27), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n600_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n310_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n257_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n616_), .B1(new_n620_), .B2(KEYINPUT17), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(KEYINPUT17), .B2(new_n616_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n620_), .A2(KEYINPUT77), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n228_), .A2(new_n303_), .A3(new_n261_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n313_), .B(KEYINPUT15), .ZN(new_n627_));
  INV_X1    g426(.A(new_n250_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n626_), .B(KEYINPUT72), .C1(new_n627_), .C2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT35), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n304_), .A2(new_n250_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n638_), .A2(KEYINPUT72), .A3(new_n626_), .A4(new_n632_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT74), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(G134gat), .ZN(new_n644_));
  INV_X1    g443(.A(G162gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT36), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n634_), .A2(new_n637_), .A3(new_n639_), .A4(KEYINPUT74), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n642_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n646_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(KEYINPUT36), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n640_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n649_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n625_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n298_), .A2(new_n326_), .A3(new_n611_), .A4(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n202_), .B1(new_n656_), .B2(new_n530_), .ZN(new_n657_));
  XOR2_X1   g456(.A(KEYINPUT75), .B(KEYINPUT37), .Z(new_n658_));
  NAND3_X1  g457(.A1(new_n649_), .A2(new_n652_), .A3(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n640_), .A2(KEYINPUT73), .A3(new_n651_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT73), .B1(new_n640_), .B2(new_n651_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n647_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n640_), .A2(new_n663_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n661_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT37), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n659_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(KEYINPUT78), .A3(new_n624_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT78), .B1(new_n667_), .B2(new_n624_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT71), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n289_), .A2(new_n290_), .A3(new_n203_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT13), .B1(new_n293_), .B2(new_n294_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n291_), .A2(new_n295_), .A3(KEYINPUT71), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT79), .B1(new_n671_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT78), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT73), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n652_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n664_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n660_), .ZN(new_n683_));
  AOI22_X1  g482(.A1(new_n653_), .A2(new_n658_), .B1(new_n683_), .B2(KEYINPUT37), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n679_), .B1(new_n684_), .B2(new_n625_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n668_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT79), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n298_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n678_), .A2(new_n326_), .A3(new_n688_), .A4(new_n611_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n530_), .A2(new_n202_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n657_), .B1(new_n691_), .B2(KEYINPUT38), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT38), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n693_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT104), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n696_), .B(new_n693_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n692_), .A2(new_n695_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT105), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n692_), .A2(new_n695_), .A3(new_n700_), .A4(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1324gat));
  NAND2_X1  g501(.A1(new_n603_), .A2(new_n609_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OR3_X1    g503(.A1(new_n689_), .A2(G8gat), .A3(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G8gat), .B1(new_n655_), .B2(new_n704_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n706_), .A2(KEYINPUT106), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(KEYINPUT106), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(KEYINPUT39), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT39), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n706_), .A2(KEYINPUT106), .A3(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n705_), .A2(new_n709_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT40), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n705_), .A2(new_n709_), .A3(KEYINPUT40), .A4(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1325gat));
  OAI21_X1  g515(.A(G15gat), .B1(new_n655_), .B2(new_n570_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT41), .Z(new_n718_));
  OR2_X1    g517(.A1(new_n570_), .A2(G15gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n689_), .B2(new_n719_), .ZN(G1326gat));
  INV_X1    g519(.A(new_n598_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G22gat), .B1(new_n655_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT42), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n721_), .A2(G22gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n689_), .B2(new_n724_), .ZN(G1327gat));
  AND4_X1   g524(.A1(new_n625_), .A2(new_n675_), .A3(new_n676_), .A4(new_n326_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n611_), .B2(new_n684_), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT43), .B(new_n667_), .C1(new_n600_), .C2(new_n610_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n726_), .B(KEYINPUT44), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n530_), .A3(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n734_), .A2(KEYINPUT107), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(KEYINPUT107), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(G29gat), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n653_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n600_), .B2(new_n610_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n726_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n530_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(G29gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n737_), .B1(new_n741_), .B2(new_n743_), .ZN(G1328gat));
  NAND3_X1  g543(.A1(new_n732_), .A2(new_n703_), .A3(new_n733_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT108), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n732_), .A2(new_n747_), .A3(new_n703_), .A4(new_n733_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(G36gat), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(G36gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n740_), .A2(new_n750_), .A3(new_n703_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT45), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n749_), .A2(KEYINPUT46), .A3(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1329gat));
  XNOR2_X1  g556(.A(KEYINPUT109), .B(G43gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n741_), .B2(new_n570_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n732_), .A2(new_n733_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n605_), .A2(G43gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n759_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g562(.A(G50gat), .B1(new_n760_), .B2(new_n721_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n740_), .A2(new_n302_), .A3(new_n598_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1331gat));
  NOR2_X1   g565(.A1(new_n298_), .A2(new_n326_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(new_n611_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n686_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n769_), .A2(new_n742_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n326_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n677_), .A2(new_n771_), .A3(new_n611_), .A4(new_n654_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n773_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n530_), .A3(new_n775_), .ZN(new_n776_));
  MUX2_X1   g575(.A(new_n770_), .B(new_n776_), .S(G57gat), .Z(G1332gat));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n703_), .A3(new_n775_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G64gat), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT111), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n781_), .A3(G64gat), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT48), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OR3_X1    g584(.A1(new_n769_), .A2(G64gat), .A3(new_n704_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n780_), .A2(KEYINPUT48), .A3(new_n782_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(G1333gat));
  NAND3_X1  g587(.A1(new_n774_), .A2(new_n571_), .A3(new_n775_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(G71gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G71gat), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n570_), .A2(G71gat), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT112), .Z(new_n794_));
  OAI22_X1  g593(.A1(new_n791_), .A2(new_n792_), .B1(new_n769_), .B2(new_n794_), .ZN(G1334gat));
  OR3_X1    g594(.A1(new_n769_), .A2(G78gat), .A3(new_n721_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n774_), .A2(new_n598_), .A3(new_n775_), .ZN(new_n797_));
  XOR2_X1   g596(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(G78gat), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G78gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT114), .B(new_n796_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1335gat));
  NAND3_X1  g604(.A1(new_n677_), .A2(new_n625_), .A3(new_n771_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n739_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n808_), .A2(G85gat), .A3(new_n742_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n767_), .A2(new_n810_), .A3(new_n625_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n806_), .A2(KEYINPUT116), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n728_), .A2(new_n729_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT115), .ZN(new_n815_));
  OR3_X1    g614(.A1(new_n728_), .A2(new_n729_), .A3(KEYINPUT115), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n813_), .A2(new_n815_), .A3(new_n816_), .A4(new_n530_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n809_), .B1(new_n817_), .B2(G85gat), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT117), .ZN(G1336gat));
  INV_X1    g618(.A(new_n808_), .ZN(new_n820_));
  AOI21_X1  g619(.A(G92gat), .B1(new_n820_), .B2(new_n703_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n813_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(new_n704_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n823_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g623(.A(G99gat), .B1(new_n822_), .B2(new_n570_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n242_), .A2(new_n244_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n820_), .A2(new_n827_), .A3(new_n605_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT51), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n825_), .A2(new_n831_), .A3(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1338gat));
  OR3_X1    g632(.A1(new_n808_), .A2(G106gat), .A3(new_n721_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n814_), .A2(new_n811_), .A3(new_n598_), .A4(new_n812_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(G106gat), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n835_), .B2(G106gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n834_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT53), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n842_), .B(new_n834_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1339gat));
  AND2_X1   g643(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n845_));
  NOR2_X1   g644(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n667_), .A2(new_n624_), .A3(new_n771_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n291_), .A2(new_n295_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n848_), .A2(new_n849_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n845_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n227_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n225_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n261_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n258_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n266_), .B2(new_n265_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n260_), .B1(new_n857_), .B2(new_n259_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n268_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n857_), .A2(KEYINPUT55), .A3(new_n260_), .A4(new_n259_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT56), .B1(new_n862_), .B2(new_n284_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864_));
  AOI211_X1 g663(.A(new_n864_), .B(new_n276_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n315_), .A2(new_n312_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n311_), .B1(new_n313_), .B2(new_n310_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n323_), .B(new_n867_), .C1(new_n868_), .C2(new_n312_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n869_), .A2(new_n325_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(KEYINPUT58), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n866_), .A2(new_n281_), .A3(new_n870_), .A4(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n281_), .B(new_n870_), .C1(new_n863_), .C2(new_n865_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n872_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n684_), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n870_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n281_), .B(new_n326_), .C1(new_n863_), .C2(new_n865_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n653_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n877_), .B1(KEYINPUT57), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(KEYINPUT57), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n881_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n850_), .B(new_n852_), .C1(new_n886_), .C2(new_n624_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n703_), .A2(new_n742_), .A3(new_n606_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G113gat), .B1(new_n889_), .B2(new_n326_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n852_), .A2(new_n850_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n881_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n884_), .A2(new_n885_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n877_), .B(KEYINPUT121), .C1(KEYINPUT57), .C2(new_n880_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n893_), .B1(new_n898_), .B2(new_n625_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n888_), .A2(new_n891_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n892_), .A2(new_n901_), .A3(new_n771_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n890_), .B1(new_n902_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g702(.A(G120gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n298_), .B2(KEYINPUT60), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n889_), .B(new_n905_), .C1(KEYINPUT60), .C2(new_n904_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n892_), .A2(new_n901_), .A3(new_n298_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n904_), .ZN(G1341gat));
  AOI21_X1  g707(.A(G127gat), .B1(new_n889_), .B2(new_n624_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n892_), .A2(new_n901_), .A3(new_n452_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n624_), .ZN(G1342gat));
  AOI21_X1  g710(.A(G134gat), .B1(new_n889_), .B2(new_n653_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n892_), .A2(new_n901_), .A3(new_n453_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n684_), .ZN(G1343gat));
  INV_X1    g713(.A(new_n604_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n703_), .A2(new_n742_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n881_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n624_), .B1(new_n917_), .B2(new_n896_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n915_), .B(new_n916_), .C1(new_n918_), .C2(new_n893_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n326_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g721(.A1(new_n919_), .A2(new_n298_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT122), .B(G148gat), .Z(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(KEYINPUT123), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n923_), .B(new_n925_), .ZN(G1345gat));
  NOR2_X1   g725(.A1(new_n919_), .A2(new_n625_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT61), .B(G155gat), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1346gat));
  NAND3_X1  g728(.A1(new_n920_), .A2(G162gat), .A3(new_n684_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n645_), .B1(new_n919_), .B2(new_n738_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT124), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(new_n934_), .A3(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n704_), .A2(new_n530_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n571_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT125), .ZN(new_n939_));
  NOR4_X1   g738(.A1(new_n899_), .A2(new_n771_), .A3(new_n598_), .A4(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n941_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n940_), .B2(new_n383_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n940_), .A2(new_n364_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n944_), .A3(new_n945_), .ZN(G1348gat));
  NOR2_X1   g745(.A1(new_n899_), .A2(new_n598_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n939_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n947_), .A2(new_n677_), .A3(new_n948_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n887_), .A2(new_n721_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n939_), .A2(new_n275_), .A3(new_n298_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n949_), .A2(new_n275_), .B1(new_n950_), .B2(new_n951_), .ZN(G1349gat));
  NAND3_X1  g751(.A1(new_n950_), .A2(new_n624_), .A3(new_n948_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n939_), .A2(new_n625_), .A3(new_n379_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n953_), .A2(new_n374_), .B1(new_n947_), .B2(new_n954_), .ZN(G1350gat));
  NAND4_X1  g754(.A1(new_n947_), .A2(new_n653_), .A3(new_n380_), .A4(new_n948_), .ZN(new_n956_));
  NOR4_X1   g755(.A1(new_n899_), .A2(new_n667_), .A3(new_n598_), .A4(new_n939_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n957_), .B2(new_n375_), .ZN(G1351gat));
  OAI211_X1 g757(.A(new_n915_), .B(new_n937_), .C1(new_n918_), .C2(new_n893_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(KEYINPUT126), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n887_), .A2(new_n961_), .A3(new_n915_), .A4(new_n937_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n960_), .A2(new_n962_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n963_), .A2(new_n326_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(G197gat), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n963_), .A2(new_n333_), .A3(new_n326_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1352gat));
  NAND2_X1  g766(.A1(new_n963_), .A2(new_n677_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n272_), .A2(KEYINPUT127), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(new_n970_));
  OAI211_X1 g769(.A(new_n963_), .B(new_n677_), .C1(KEYINPUT127), .C2(new_n272_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(G1353gat));
  NOR2_X1   g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  AND2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  OAI211_X1 g773(.A(new_n963_), .B(new_n624_), .C1(new_n973_), .C2(new_n974_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n625_), .B1(new_n960_), .B2(new_n962_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n975_), .B1(new_n976_), .B2(new_n973_), .ZN(G1354gat));
  AOI21_X1  g776(.A(G218gat), .B1(new_n963_), .B2(new_n653_), .ZN(new_n978_));
  INV_X1    g777(.A(G218gat), .ZN(new_n979_));
  AOI211_X1 g778(.A(new_n979_), .B(new_n667_), .C1(new_n960_), .C2(new_n962_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n978_), .A2(new_n980_), .ZN(G1355gat));
endmodule


