//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n204_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT77), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT23), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  OR3_X1    g017(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n204_), .A2(new_n209_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(KEYINPUT77), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n212_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n217_), .A2(new_n224_), .ZN(new_n225_));
  OAI221_X1 g024(.A(new_n225_), .B1(G183gat), .B2(G190gat), .C1(new_n218_), .C2(KEYINPUT78), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(G169gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G43gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n230_), .B(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n233_), .B(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  INV_X1    g037(.A(G15gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT30), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT31), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n237_), .B(new_n242_), .Z(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(G155gat), .B(G162gat), .Z(new_n246_));
  INV_X1    g045(.A(G141gat), .ZN(new_n247_));
  INV_X1    g046(.A(G148gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT2), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G141gat), .A2(G148gat), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n249_), .A2(KEYINPUT3), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(KEYINPUT3), .B2(new_n249_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT79), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n246_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n246_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n249_), .A4(new_n251_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(KEYINPUT88), .A3(new_n236_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n262_), .B(KEYINPUT4), .C1(new_n236_), .C2(new_n261_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n261_), .A2(KEYINPUT88), .A3(new_n264_), .A4(new_n236_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n245_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n261_), .B(new_n236_), .Z(new_n268_));
  INV_X1    g067(.A(new_n245_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G1gat), .B(G29gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G85gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT0), .B(G57gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n267_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(new_n266_), .B2(new_n270_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT90), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n267_), .A2(new_n271_), .A3(KEYINPUT90), .A4(new_n276_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n244_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n286_));
  NOR2_X1   g085(.A1(new_n261_), .A2(KEYINPUT29), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT80), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n287_), .A2(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n286_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n291_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n286_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G228gat), .A2(G233gat), .ZN(new_n297_));
  INV_X1    g096(.A(G78gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G106gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n292_), .A2(new_n295_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT83), .ZN(new_n306_));
  INV_X1    g105(.A(G204gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(G197gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(G197gat), .ZN(new_n309_));
  INV_X1    g108(.A(G197gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(KEYINPUT83), .A3(G204gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n312_), .A2(KEYINPUT21), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT21), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(G204gat), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(new_n309_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT82), .Z(new_n319_));
  NOR2_X1   g118(.A1(new_n314_), .A2(new_n316_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n315_), .A2(new_n319_), .B1(new_n312_), .B2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(KEYINPUT29), .B2(new_n261_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G22gat), .B(G50gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n305_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n302_), .A2(new_n324_), .A3(new_n304_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n225_), .B(new_n219_), .C1(new_n218_), .C2(KEYINPUT78), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT85), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n210_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n218_), .B1(G183gat), .B2(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n338_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n228_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n321_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n315_), .A2(new_n319_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n320_), .A2(new_n312_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT20), .B1(new_n345_), .B2(new_n230_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n333_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G8gat), .B(G36gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n345_), .B2(new_n230_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n336_), .A2(new_n321_), .A3(new_n341_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n356_), .A3(new_n332_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n347_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n347_), .B2(new_n357_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n329_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT91), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n342_), .A2(new_n346_), .A3(new_n333_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n332_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n352_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT27), .A3(new_n358_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n361_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n362_), .B1(new_n361_), .B2(new_n366_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n328_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT92), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n361_), .A2(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT91), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n361_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT92), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n328_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n285_), .B1(new_n370_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT33), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n278_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT89), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n359_), .A2(new_n360_), .ZN(new_n381_));
  OAI211_X1 g180(.A(KEYINPUT33), .B(new_n275_), .C1(new_n266_), .C2(new_n270_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n263_), .A2(new_n245_), .A3(new_n265_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n268_), .A2(new_n269_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(new_n276_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(KEYINPUT32), .B(new_n353_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n347_), .A2(new_n388_), .A3(new_n357_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  OAI22_X1  g189(.A1(new_n380_), .A2(new_n386_), .B1(new_n282_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n328_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n326_), .A2(new_n327_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n393_), .A2(new_n282_), .A3(new_n361_), .A4(new_n366_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n243_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n377_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G8gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT75), .ZN(new_n398_));
  INV_X1    g197(.A(G22gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n239_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G15gat), .A2(G22gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G1gat), .A2(G8gat), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n400_), .A2(new_n401_), .B1(KEYINPUT14), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n398_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G29gat), .B(G36gat), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(KEYINPUT74), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(KEYINPUT74), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G43gat), .B(G50gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n404_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G229gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n404_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT15), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n411_), .A2(KEYINPUT15), .A3(new_n412_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n416_), .B1(new_n404_), .B2(new_n413_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n414_), .A2(new_n416_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G141gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G169gat), .B(G197gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n424_), .B(new_n425_), .Z(new_n426_));
  OR2_X1    g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n423_), .A2(new_n426_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n396_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G230gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT64), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT9), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(G85gat), .A3(G92gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G85gat), .B(G92gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n435_), .B1(new_n436_), .B2(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT66), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT66), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n439_), .B(new_n435_), .C1(new_n436_), .C2(new_n434_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT10), .B(G99gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT65), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n441_), .B(new_n445_), .C1(G106gat), .C2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT8), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT69), .ZN(new_n450_));
  INV_X1    g249(.A(G99gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n300_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n453_));
  OR2_X1    g252(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n450_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n456_), .B1(new_n460_), .B2(new_n457_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n454_), .A2(new_n452_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT69), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n463_), .A3(new_n445_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n436_), .B(KEYINPUT68), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n449_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n462_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(new_n444_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT68), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n436_), .B(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n468_), .A2(new_n470_), .A3(KEYINPUT8), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n448_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G57gat), .B(G64gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n473_), .A2(KEYINPUT11), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT70), .B(G71gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n475_), .A2(G78gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(G78gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n474_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n473_), .B(KEYINPUT11), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n476_), .A2(new_n477_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n472_), .A2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n448_), .B(new_n481_), .C1(new_n466_), .C2(new_n471_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n433_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT12), .B1(new_n472_), .B2(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n484_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(KEYINPUT12), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n485_), .B1(new_n488_), .B2(new_n433_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G120gat), .B(G148gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT5), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(KEYINPUT71), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT72), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n489_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n489_), .A2(new_n496_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT13), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(KEYINPUT13), .A3(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n472_), .A2(new_n420_), .A3(new_n419_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n465_), .B(new_n449_), .C1(new_n467_), .C2(new_n444_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n444_), .B1(new_n467_), .B2(new_n450_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n470_), .B1(new_n507_), .B2(new_n463_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n508_), .B2(new_n449_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n413_), .A3(new_n448_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n505_), .B(new_n510_), .C1(KEYINPUT35), .C2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(KEYINPUT35), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G190gat), .B(G218gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G134gat), .B(G162gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT36), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n519_), .A2(KEYINPUT36), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n516_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n516_), .A2(new_n520_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT37), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n481_), .B(new_n528_), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n404_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G127gat), .B(G155gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G183gat), .B(G211gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n535_), .A2(KEYINPUT17), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n535_), .B(KEYINPUT17), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n530_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n527_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n431_), .A2(new_n504_), .A3(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT93), .Z(new_n544_));
  INV_X1    g343(.A(G1gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n283_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n548_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n396_), .A2(new_n524_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n503_), .A2(new_n430_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n540_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT95), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(G1gat), .B1(new_n555_), .B2(new_n282_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n549_), .A2(new_n550_), .A3(new_n556_), .ZN(G1324gat));
  INV_X1    g356(.A(G8gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n374_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n544_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT39), .ZN(new_n561_));
  INV_X1    g360(.A(new_n555_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n559_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n563_), .B2(G8gat), .ZN(new_n564_));
  AOI211_X1 g363(.A(KEYINPUT39), .B(new_n558_), .C1(new_n562_), .C2(new_n559_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n560_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g366(.A(new_n543_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n569_));
  OAI21_X1  g368(.A(G15gat), .B1(new_n555_), .B2(new_n244_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT41), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(new_n571_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n569_), .B1(new_n572_), .B2(new_n573_), .ZN(G1326gat));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n399_), .A3(new_n393_), .ZN(new_n575_));
  OAI21_X1  g374(.A(G22gat), .B1(new_n555_), .B2(new_n328_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n576_), .A2(KEYINPUT42), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(KEYINPUT42), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n575_), .B1(new_n577_), .B2(new_n578_), .ZN(G1327gat));
  NAND2_X1  g378(.A1(new_n524_), .A2(new_n541_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT97), .Z(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n503_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n431_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(G29gat), .B1(new_n584_), .B2(new_n283_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n527_), .B1(new_n377_), .B2(new_n395_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT43), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT43), .B(new_n527_), .C1(new_n377_), .C2(new_n395_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n541_), .A3(new_n552_), .A4(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT44), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n540_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n593_), .A2(KEYINPUT96), .A3(new_n552_), .A4(new_n589_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n590_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n592_), .A2(new_n594_), .B1(KEYINPUT44), .B2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n283_), .A2(G29gat), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n585_), .B1(new_n596_), .B2(new_n597_), .ZN(G1328gat));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT99), .B(KEYINPUT45), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n374_), .A2(G36gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OR3_X1    g401(.A1(new_n583_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n583_), .B2(new_n602_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(G36gat), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT44), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n559_), .B1(new_n590_), .B2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n594_), .B2(new_n592_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n606_), .B1(new_n609_), .B2(KEYINPUT98), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n592_), .A2(new_n594_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n605_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT100), .B(KEYINPUT46), .Z(new_n617_));
  OAI21_X1  g416(.A(new_n599_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(KEYINPUT46), .ZN(new_n619_));
  INV_X1    g418(.A(new_n605_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n611_), .A2(new_n612_), .A3(KEYINPUT98), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(G36gat), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n609_), .A2(KEYINPUT98), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n620_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n617_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(KEYINPUT101), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n618_), .A2(new_n619_), .A3(new_n626_), .ZN(G1329gat));
  NOR3_X1   g426(.A1(new_n583_), .A2(G43gat), .A3(new_n244_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n596_), .A2(new_n243_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n629_), .B2(G43gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n630_), .B(new_n631_), .Z(G1330gat));
  OR3_X1    g431(.A1(new_n583_), .A2(G50gat), .A3(new_n328_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n596_), .A2(new_n393_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(KEYINPUT103), .ZN(new_n635_));
  OAI21_X1  g434(.A(G50gat), .B1(new_n634_), .B2(KEYINPUT103), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n633_), .B1(new_n635_), .B2(new_n636_), .ZN(G1331gat));
  NAND2_X1  g436(.A1(new_n542_), .A2(new_n503_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT104), .Z(new_n639_));
  NOR2_X1   g438(.A1(new_n396_), .A2(new_n429_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G57gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(new_n283_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n540_), .A2(new_n430_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n504_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n551_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G57gat), .B1(new_n647_), .B2(new_n282_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(G1332gat));
  INV_X1    g448(.A(G64gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n642_), .A2(new_n650_), .A3(new_n559_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G64gat), .B1(new_n647_), .B2(new_n374_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT48), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1333gat));
  INV_X1    g453(.A(G71gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n642_), .A2(new_n655_), .A3(new_n243_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n647_), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT49), .B(new_n655_), .C1(new_n657_), .C2(new_n243_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT49), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n243_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(G71gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n656_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT105), .Z(G1334gat));
  NAND3_X1  g462(.A1(new_n642_), .A2(new_n298_), .A3(new_n393_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G78gat), .B1(new_n647_), .B2(new_n328_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT50), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1335gat));
  NOR3_X1   g466(.A1(new_n641_), .A2(new_n504_), .A3(new_n581_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n282_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n593_), .A2(new_n430_), .A3(new_n503_), .A4(new_n589_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n283_), .A2(G85gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT106), .ZN(new_n673_));
  OAI22_X1  g472(.A1(new_n670_), .A2(G85gat), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT107), .ZN(G1336gat));
  OAI21_X1  g474(.A(G92gat), .B1(new_n671_), .B2(new_n374_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n374_), .A2(G92gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n669_), .B2(new_n677_), .ZN(G1337gat));
  INV_X1    g477(.A(KEYINPUT51), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(KEYINPUT108), .ZN(new_n680_));
  INV_X1    g479(.A(new_n671_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n451_), .B1(new_n681_), .B2(new_n243_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n244_), .A2(new_n447_), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n680_), .B(new_n682_), .C1(new_n668_), .C2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n679_), .A2(KEYINPUT108), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n684_), .B(new_n685_), .Z(G1338gat));
  OAI21_X1  g485(.A(G106gat), .B1(new_n671_), .B2(new_n328_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(KEYINPUT52), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(KEYINPUT52), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n668_), .A2(new_n300_), .A3(new_n393_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1339gat));
  INV_X1    g493(.A(G113gat), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n370_), .A2(new_n376_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n283_), .A2(new_n243_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT119), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(KEYINPUT116), .B2(KEYINPUT57), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n414_), .A2(new_n415_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n415_), .B1(new_n404_), .B2(new_n413_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n421_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n426_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT115), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT115), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n704_), .A2(new_n706_), .A3(new_n710_), .A4(new_n707_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(new_n428_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT12), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n716_), .B2(new_n486_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n433_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n484_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n481_), .B1(new_n509_), .B2(new_n448_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT12), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n472_), .A2(new_n482_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n715_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n721_), .A2(KEYINPUT112), .A3(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n717_), .A2(new_n718_), .A3(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n721_), .A2(KEYINPUT55), .A3(new_n433_), .A4(new_n723_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n488_), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n433_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n721_), .A2(new_n433_), .A3(new_n723_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n725_), .A2(new_n728_), .A3(new_n729_), .A4(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT114), .B1(new_n733_), .B2(new_n493_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT56), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n733_), .B2(new_n493_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n489_), .A2(new_n494_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n429_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n734_), .A2(new_n736_), .A3(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n733_), .A2(KEYINPUT114), .A3(new_n735_), .A4(new_n493_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n713_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n522_), .A2(new_n523_), .B1(new_n701_), .B2(KEYINPUT57), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n703_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n734_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n733_), .A2(new_n493_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT56), .ZN(new_n746_));
  INV_X1    g545(.A(new_n738_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n744_), .A2(new_n746_), .A3(new_n740_), .A4(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n713_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n742_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n702_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n743_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n733_), .A2(new_n735_), .A3(new_n493_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n712_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT117), .B(KEYINPUT58), .C1(new_n756_), .C2(new_n736_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n746_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT58), .B1(new_n759_), .B2(KEYINPUT117), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n527_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n753_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n541_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n645_), .B(KEYINPUT110), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n526_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n766_), .A2(KEYINPUT111), .A3(KEYINPUT54), .A4(new_n504_), .ZN(new_n767_));
  OR2_X1    g566(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n768_));
  NAND2_X1  g567(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n768_), .B(new_n769_), .C1(new_n765_), .C2(new_n503_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT59), .B(new_n700_), .C1(new_n763_), .C2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n761_), .A2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n527_), .B(KEYINPUT118), .C1(new_n758_), .C2(new_n760_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n753_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n771_), .B1(new_n777_), .B2(new_n541_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT59), .B1(new_n778_), .B2(new_n700_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT120), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n778_), .C2(new_n700_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n773_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n695_), .B1(new_n783_), .B2(new_n429_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n778_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n699_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n429_), .A2(new_n695_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT121), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n790_));
  INV_X1    g589(.A(new_n788_), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n430_), .B(new_n773_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n790_), .B(new_n791_), .C1(new_n792_), .C2(new_n695_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(G1340gat));
  INV_X1    g593(.A(new_n786_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT60), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT122), .B1(new_n796_), .B2(G120gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(G120gat), .B1(new_n503_), .B2(new_n796_), .ZN(new_n798_));
  MUX2_X1   g597(.A(new_n797_), .B(KEYINPUT122), .S(new_n798_), .Z(new_n799_));
  NAND2_X1  g598(.A1(new_n795_), .A2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n783_), .A2(new_n503_), .ZN(new_n801_));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(G1341gat));
  AOI21_X1  g602(.A(G127gat), .B1(new_n795_), .B2(new_n540_), .ZN(new_n804_));
  XOR2_X1   g603(.A(KEYINPUT123), .B(G127gat), .Z(new_n805_));
  NAND2_X1  g604(.A1(new_n540_), .A2(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT124), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n804_), .B1(new_n783_), .B2(new_n807_), .ZN(G1342gat));
  INV_X1    g607(.A(KEYINPUT125), .ZN(new_n809_));
  INV_X1    g608(.A(G134gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n783_), .B2(new_n527_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n524_), .A2(new_n810_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n786_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n813_), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n526_), .B(new_n773_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT125), .B(new_n815_), .C1(new_n816_), .C2(new_n810_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(G1343gat));
  NOR2_X1   g617(.A1(new_n328_), .A2(new_n243_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(new_n374_), .A3(new_n283_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n785_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT126), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n822_), .A2(new_n823_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n429_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g627(.A(new_n503_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g629(.A(new_n540_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT61), .B(G155gat), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1346gat));
  INV_X1    g632(.A(G162gat), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n524_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n826_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n526_), .B1(new_n836_), .B2(new_n824_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n837_), .B2(new_n834_), .ZN(G1347gat));
  NAND2_X1  g637(.A1(new_n763_), .A2(new_n772_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n285_), .A2(new_n374_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n393_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n429_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT62), .B1(new_n845_), .B2(KEYINPUT22), .ZN(new_n846_));
  OAI21_X1  g645(.A(G169gat), .B1(new_n845_), .B2(KEYINPUT62), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n207_), .B2(new_n846_), .ZN(G1348gat));
  AOI21_X1  g648(.A(G176gat), .B1(new_n844_), .B2(new_n503_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n778_), .A2(new_n393_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n841_), .A2(new_n504_), .A3(new_n208_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(G1349gat));
  NOR3_X1   g652(.A1(new_n843_), .A2(new_n202_), .A3(new_n541_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n540_), .A3(new_n840_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n213_), .B2(new_n855_), .ZN(G1350gat));
  OAI21_X1  g655(.A(G190gat), .B1(new_n843_), .B2(new_n526_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n524_), .A2(new_n203_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n843_), .B2(new_n858_), .ZN(G1351gat));
  AND4_X1   g658(.A1(new_n282_), .A2(new_n785_), .A3(new_n559_), .A4(new_n819_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n429_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n503_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g663(.A(KEYINPUT63), .B(G211gat), .C1(new_n860_), .C2(new_n540_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n860_), .A2(new_n540_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT63), .B(G211gat), .Z(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(G1354gat));
  NAND2_X1  g667(.A1(new_n860_), .A2(new_n524_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT127), .B(G218gat), .Z(new_n870_));
  NOR2_X1   g669(.A1(new_n526_), .A2(new_n870_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n869_), .A2(new_n870_), .B1(new_n860_), .B2(new_n871_), .ZN(G1355gat));
endmodule


