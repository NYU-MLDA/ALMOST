//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT20), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT84), .B(G204gat), .ZN(new_n207_));
  INV_X1    g006(.A(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI22_X1  g008(.A1(new_n209_), .A2(KEYINPUT85), .B1(new_n208_), .B2(G204gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(KEYINPUT85), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT21), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G197gat), .A2(G204gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n213_), .B1(new_n207_), .B2(G197gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT21), .ZN(new_n215_));
  XOR2_X1   g014(.A(G211gat), .B(G218gat), .Z(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(KEYINPUT21), .A3(new_n216_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT75), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226_));
  INV_X1    g025(.A(G169gat), .ZN(new_n227_));
  INV_X1    g026(.A(G176gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n225_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(new_n226_), .B2(new_n225_), .ZN(new_n231_));
  INV_X1    g030(.A(G183gat), .ZN(new_n232_));
  INV_X1    g031(.A(G190gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT23), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT76), .ZN(new_n235_));
  OR3_X1    g034(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT23), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT26), .B(G190gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT74), .B1(new_n232_), .B2(KEYINPUT25), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT25), .B(G183gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n238_), .B(new_n239_), .C1(new_n240_), .C2(KEYINPUT74), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n231_), .A2(new_n237_), .A3(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT22), .B(G169gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n228_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT77), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n236_), .A2(new_n234_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n232_), .A2(new_n233_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n229_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n206_), .B1(new_n220_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n237_), .A2(new_n248_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n253_), .B(new_n244_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n240_), .A2(new_n238_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n231_), .A2(new_n247_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(new_n220_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(KEYINPUT88), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(KEYINPUT88), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n205_), .B(new_n252_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT90), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n220_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n268_), .B(KEYINPUT20), .C1(new_n251_), .C2(new_n220_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n204_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n261_), .A2(new_n267_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n267_), .B1(new_n261_), .B2(new_n270_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n202_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G141gat), .A2(G148gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT80), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT2), .ZN(new_n281_));
  OR3_X1    g080(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  INV_X1    g081(.A(G141gat), .ZN(new_n283_));
  INV_X1    g082(.A(G148gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT3), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n281_), .A2(new_n282_), .A3(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n280_), .A2(KEYINPUT2), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n278_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n275_), .A2(KEYINPUT1), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n275_), .B1(new_n277_), .B2(KEYINPUT1), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT79), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(new_n294_), .B2(new_n293_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n279_), .A3(new_n285_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n291_), .A2(KEYINPUT82), .A3(new_n297_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G127gat), .B(G134gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G120gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(new_n298_), .B2(new_n304_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT4), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n307_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(G85gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT0), .B(G57gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n306_), .A2(new_n308_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n312_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n318_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n316_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT92), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n220_), .B1(new_n257_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n322_), .B2(new_n257_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n205_), .B1(new_n324_), .B2(new_n252_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n269_), .A2(new_n204_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n271_), .B(KEYINPUT27), .C1(new_n327_), .C2(new_n267_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n274_), .A2(new_n319_), .A3(new_n321_), .A4(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G71gat), .B(G99gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G43gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(G15gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n331_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n251_), .B(KEYINPUT30), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n336_), .A2(new_n337_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n338_), .B2(new_n335_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n304_), .B(KEYINPUT31), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G22gat), .B(G50gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n220_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(KEYINPUT86), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(KEYINPUT86), .B2(new_n347_), .ZN(new_n349_));
  INV_X1    g148(.A(G228gat), .ZN(new_n350_));
  OR2_X1    g149(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n346_), .A2(new_n353_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n300_), .A2(new_n301_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n345_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n358_), .A3(new_n345_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G78gat), .B(G106gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n362_), .B(KEYINPUT87), .Z(new_n363_));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n356_), .A2(new_n364_), .A3(new_n357_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n363_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n363_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(new_n365_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n360_), .A2(new_n361_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n361_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n371_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n359_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n343_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n342_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n341_), .B(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n360_), .A2(new_n368_), .A3(new_n371_), .A4(new_n361_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n374_), .B1(new_n373_), .B2(new_n359_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n329_), .B1(new_n376_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n321_), .A2(new_n319_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n261_), .A2(new_n270_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n267_), .A2(KEYINPUT32), .ZN(new_n385_));
  MUX2_X1   g184(.A(new_n327_), .B(new_n384_), .S(new_n385_), .Z(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT93), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n317_), .B1(new_n312_), .B2(new_n318_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n389_), .A2(KEYINPUT33), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(KEYINPUT33), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n309_), .B1(new_n307_), .B2(new_n311_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n317_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(KEYINPUT91), .B2(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n393_), .A2(KEYINPUT91), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n272_), .A2(new_n273_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n390_), .A2(new_n391_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT93), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n383_), .A2(new_n399_), .A3(new_n386_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n388_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n372_), .A2(new_n375_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(new_n378_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n382_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G113gat), .B(G141gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G169gat), .B(G197gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G229gat), .A2(G233gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G15gat), .B(G22gat), .ZN(new_n411_));
  INV_X1    g210(.A(G1gat), .ZN(new_n412_));
  INV_X1    g211(.A(G8gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT14), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G1gat), .B(G8gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G29gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G43gat), .B(G50gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n417_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT73), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n422_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n410_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n418_), .B(new_n419_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT15), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n417_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n417_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n426_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n430_), .A3(new_n410_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n409_), .B1(new_n425_), .B2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n421_), .B(KEYINPUT73), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n431_), .B(new_n408_), .C1(new_n434_), .C2(new_n410_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n405_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G231gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n417_), .B(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(G71gat), .A2(G78gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G71gat), .A2(G78gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G57gat), .B(G64gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(KEYINPUT11), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT65), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n444_), .B2(KEYINPUT11), .ZN(new_n447_));
  INV_X1    g246(.A(G64gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G57gat), .ZN(new_n449_));
  INV_X1    g248(.A(G57gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G64gat), .ZN(new_n451_));
  AND4_X1   g250(.A1(new_n446_), .A2(new_n449_), .A3(new_n451_), .A4(KEYINPUT11), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n445_), .B1(new_n447_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n451_), .A3(KEYINPUT11), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT65), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(new_n451_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT11), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n449_), .A2(new_n451_), .A3(new_n446_), .A4(KEYINPUT11), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n455_), .A2(new_n458_), .A3(new_n443_), .A4(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n453_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n440_), .B(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G127gat), .B(G155gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G183gat), .B(G211gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT17), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n467_), .A2(KEYINPUT17), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n462_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n462_), .A2(new_n468_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n472_), .B(KEYINPUT71), .Z(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT10), .B(G99gat), .Z(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n477_), .A2(KEYINPUT9), .ZN(new_n478_));
  AND3_X1   g277(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(G85gat), .A2(G92gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(KEYINPUT9), .A3(new_n477_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n476_), .A2(new_n478_), .A3(new_n481_), .A4(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(G99gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n475_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT64), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n485_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n488_), .A2(new_n481_), .A3(new_n489_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT8), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n482_), .A2(new_n477_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n493_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n484_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G232gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT34), .ZN(new_n501_));
  OAI22_X1  g300(.A1(new_n499_), .A2(new_n420_), .B1(KEYINPUT35), .B2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n499_), .A2(new_n427_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(KEYINPUT35), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n504_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G190gat), .B(G218gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G134gat), .B(G162gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT36), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n510_), .B(KEYINPUT36), .Z(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n507_), .B2(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT37), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(KEYINPUT37), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n473_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G120gat), .B(G148gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G176gat), .B(G204gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G230gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  AND4_X1   g324(.A1(new_n476_), .A2(new_n478_), .A3(new_n481_), .A4(new_n483_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n489_), .ZN(new_n531_));
  NOR4_X1   g330(.A1(KEYINPUT64), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n491_), .B1(new_n490_), .B2(new_n485_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT8), .B1(new_n534_), .B2(new_n495_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n493_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n526_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n525_), .B1(new_n537_), .B2(new_n461_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n461_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n499_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n524_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n499_), .A2(new_n525_), .A3(new_n539_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n461_), .B(new_n484_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n524_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n544_), .B2(new_n524_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n537_), .A2(KEYINPUT12), .A3(new_n461_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n499_), .B2(new_n539_), .ZN(new_n550_));
  OAI22_X1  g349(.A1(new_n546_), .A2(new_n547_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n523_), .B1(new_n552_), .B2(KEYINPUT68), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(KEYINPUT68), .B2(new_n552_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n552_), .B2(new_n522_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n544_), .A2(new_n524_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT67), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n544_), .A2(new_n545_), .A3(new_n524_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT12), .B1(new_n537_), .B2(new_n461_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n499_), .A2(new_n549_), .A3(new_n539_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n560_), .A2(new_n563_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(KEYINPUT69), .A3(new_n523_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n556_), .A2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n554_), .A2(KEYINPUT13), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT13), .B1(new_n554_), .B2(new_n566_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n518_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT72), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n438_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n412_), .A3(new_n383_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT38), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n515_), .A2(KEYINPUT95), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n512_), .B(new_n577_), .C1(new_n507_), .C2(new_n514_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n405_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n581_));
  INV_X1    g380(.A(new_n569_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n581_), .B1(new_n582_), .B2(new_n437_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n472_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n569_), .A2(KEYINPUT94), .A3(new_n436_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n580_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n383_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G1gat), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n573_), .A2(new_n574_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n575_), .A2(new_n590_), .A3(new_n591_), .ZN(G1324gat));
  NAND2_X1  g391(.A1(new_n274_), .A2(new_n328_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n572_), .A2(new_n413_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n587_), .A2(new_n593_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n596_), .B2(G8gat), .ZN(new_n597_));
  AOI211_X1 g396(.A(KEYINPUT39), .B(new_n413_), .C1(new_n587_), .C2(new_n593_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT40), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(G1325gat));
  NAND3_X1  g400(.A1(new_n572_), .A2(new_n333_), .A3(new_n378_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G15gat), .B1(new_n588_), .B2(new_n343_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT41), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n603_), .A2(new_n604_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(G1326gat));
  INV_X1    g406(.A(G22gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n572_), .A2(new_n608_), .A3(new_n403_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G22gat), .B1(new_n588_), .B2(new_n402_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(KEYINPUT42), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(KEYINPUT42), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(G1327gat));
  NAND2_X1  g412(.A1(new_n401_), .A2(new_n404_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n382_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n473_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n579_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n582_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n436_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT98), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n438_), .A2(new_n622_), .A3(new_n619_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(G29gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n383_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT99), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n583_), .A2(new_n473_), .A3(new_n585_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n516_), .A2(new_n517_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT43), .B1(new_n631_), .B2(KEYINPUT96), .ZN(new_n632_));
  INV_X1    g431(.A(new_n631_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n616_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n632_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n405_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n630_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n616_), .A2(new_n633_), .A3(new_n632_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n635_), .B1(new_n405_), .B2(new_n631_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n629_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT97), .B1(new_n643_), .B2(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT44), .B(new_n630_), .C1(new_n634_), .C2(new_n636_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(new_n383_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n628_), .B1(new_n647_), .B2(new_n625_), .ZN(G1328gat));
  INV_X1    g447(.A(new_n593_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(G36gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n621_), .A2(new_n623_), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT45), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n646_), .A2(new_n593_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n644_), .B2(new_n640_), .ZN(new_n654_));
  INV_X1    g453(.A(G36gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n652_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n652_), .B(KEYINPUT46), .C1(new_n654_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1329gat));
  AND3_X1   g459(.A1(new_n646_), .A2(G43gat), .A3(new_n378_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n645_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G43gat), .B1(new_n624_), .B2(new_n378_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT47), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n645_), .B2(new_n661_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(G1330gat));
  INV_X1    g467(.A(G50gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n624_), .A2(new_n669_), .A3(new_n403_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n646_), .A2(new_n403_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n644_), .B2(new_n640_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT100), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G50gat), .B1(new_n672_), .B2(KEYINPUT100), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n670_), .B1(new_n674_), .B2(new_n675_), .ZN(G1331gat));
  NOR2_X1   g475(.A1(new_n569_), .A2(new_n436_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n617_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n580_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G57gat), .B1(new_n680_), .B2(new_n589_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n616_), .A2(new_n518_), .A3(new_n677_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n683_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n383_), .A2(new_n450_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n681_), .B1(new_n686_), .B2(new_n687_), .ZN(G1332gat));
  INV_X1    g487(.A(new_n686_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n448_), .A3(new_n593_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G64gat), .B1(new_n680_), .B2(new_n649_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT48), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1333gat));
  OAI21_X1  g492(.A(G71gat), .B1(new_n680_), .B2(new_n343_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT49), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n343_), .A2(G71gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n686_), .B2(new_n696_), .ZN(G1334gat));
  OR3_X1    g496(.A1(new_n686_), .A2(G78gat), .A3(new_n402_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n580_), .A2(new_n403_), .A3(new_n679_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G78gat), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT50), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT102), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n704_), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1335gat));
  NOR2_X1   g505(.A1(new_n617_), .A2(new_n618_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n616_), .A2(new_n707_), .A3(new_n677_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT103), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n616_), .A2(new_n710_), .A3(new_n707_), .A4(new_n677_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G85gat), .B1(new_n712_), .B2(new_n383_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n677_), .A2(new_n473_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n383_), .A2(G85gat), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT104), .Z(new_n717_));
  AOI21_X1  g516(.A(new_n713_), .B1(new_n715_), .B2(new_n717_), .ZN(G1336gat));
  INV_X1    g517(.A(G92gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n712_), .A2(new_n719_), .A3(new_n593_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n715_), .A2(new_n593_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n719_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT105), .Z(G1337gat));
  NAND3_X1  g522(.A1(new_n712_), .A2(new_n378_), .A3(new_n474_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n715_), .A2(new_n378_), .ZN(new_n726_));
  OAI221_X1 g525(.A(new_n724_), .B1(KEYINPUT106), .B2(new_n725_), .C1(new_n726_), .C2(new_n486_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(KEYINPUT106), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(G1338gat));
  XNOR2_X1  g528(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n475_), .B1(new_n715_), .B2(new_n403_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n732_), .A2(KEYINPUT52), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(KEYINPUT52), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n402_), .A2(G106gat), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n712_), .A2(KEYINPUT107), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT107), .B1(new_n712_), .B2(new_n736_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n731_), .B1(new_n735_), .B2(new_n739_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n737_), .A2(new_n738_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n741_), .A2(new_n733_), .A3(new_n734_), .A4(new_n730_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1339gat));
  NAND3_X1  g542(.A1(new_n518_), .A2(new_n437_), .A3(new_n569_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n744_), .A2(KEYINPUT109), .A3(KEYINPUT54), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(KEYINPUT54), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT109), .B1(new_n744_), .B2(KEYINPUT54), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n744_), .A2(KEYINPUT110), .A3(KEYINPUT54), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n745_), .A2(new_n748_), .A3(new_n749_), .A4(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n410_), .B1(new_n429_), .B2(new_n426_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n408_), .B1(new_n428_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n410_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n434_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n435_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n556_), .B2(new_n565_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n758_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT56), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n524_), .B1(new_n563_), .B2(new_n544_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n551_), .A2(KEYINPUT55), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n563_), .B(new_n764_), .C1(new_n547_), .C2(new_n546_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n762_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n761_), .B1(new_n766_), .B2(new_n523_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n523_), .A2(new_n761_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n766_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n759_), .A2(new_n760_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(KEYINPUT115), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(KEYINPUT115), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n759_), .A2(new_n760_), .A3(new_n774_), .A4(new_n770_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n633_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  INV_X1    g576(.A(new_n762_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n765_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n764_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(KEYINPUT112), .A3(new_n768_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n766_), .B2(new_n769_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n767_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT69), .B1(new_n564_), .B2(new_n523_), .ZN(new_n786_));
  AND4_X1   g585(.A1(KEYINPUT69), .A2(new_n543_), .A3(new_n551_), .A4(new_n523_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n436_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n566_), .A2(KEYINPUT111), .A3(new_n436_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n554_), .A2(new_n566_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n756_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n579_), .B1(new_n792_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n777_), .B1(new_n796_), .B2(KEYINPUT113), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n798_), .B(new_n579_), .C1(new_n792_), .C2(new_n795_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n776_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n796_), .A2(KEYINPUT57), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n472_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n751_), .A2(new_n802_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n381_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT59), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n801_), .B1(new_n800_), .B2(KEYINPUT116), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(new_n776_), .C1(new_n797_), .C2(new_n799_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n617_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n751_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n807_), .B(new_n804_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n806_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(G113gat), .B1(new_n814_), .B2(new_n437_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n437_), .A2(G113gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n805_), .B2(new_n816_), .ZN(G1340gat));
  INV_X1    g616(.A(G120gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n569_), .B2(KEYINPUT60), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(KEYINPUT60), .B2(new_n818_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n805_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT117), .ZN(new_n822_));
  OAI21_X1  g621(.A(G120gat), .B1(new_n814_), .B2(new_n569_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1341gat));
  INV_X1    g623(.A(G127gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n805_), .B2(new_n473_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n826_), .A2(new_n827_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n814_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n472_), .A2(new_n825_), .ZN(new_n831_));
  AOI211_X1 g630(.A(new_n828_), .B(new_n829_), .C1(new_n830_), .C2(new_n831_), .ZN(G1342gat));
  INV_X1    g631(.A(new_n805_), .ZN(new_n833_));
  AOI21_X1  g632(.A(G134gat), .B1(new_n833_), .B2(new_n579_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n633_), .A2(G134gat), .ZN(new_n835_));
  XOR2_X1   g634(.A(new_n835_), .B(KEYINPUT119), .Z(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n830_), .B2(new_n836_), .ZN(G1343gat));
  NOR3_X1   g636(.A1(new_n376_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(KEYINPUT120), .Z(new_n839_));
  NAND2_X1  g638(.A1(new_n803_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n437_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n283_), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n569_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n284_), .ZN(G1345gat));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845_));
  INV_X1    g644(.A(new_n840_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n617_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n840_), .A2(KEYINPUT121), .A3(new_n473_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT61), .B(G155gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1346gat));
  AOI21_X1  g650(.A(G162gat), .B1(new_n846_), .B2(new_n579_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n633_), .A2(G162gat), .ZN(new_n853_));
  XOR2_X1   g652(.A(new_n853_), .B(KEYINPUT122), .Z(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n846_), .B2(new_n854_), .ZN(G1347gat));
  NAND3_X1  g654(.A1(new_n593_), .A2(new_n589_), .A3(new_n378_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n403_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n436_), .B(new_n857_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n243_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(G169gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT123), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n860_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n861_), .A2(KEYINPUT123), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(KEYINPUT62), .A3(new_n862_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1348gat));
  OAI21_X1  g667(.A(new_n857_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n228_), .B1(new_n869_), .B2(new_n569_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n403_), .B1(new_n751_), .B2(new_n802_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n856_), .A2(new_n228_), .A3(new_n569_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT124), .ZN(G1349gat));
  NOR3_X1   g674(.A1(new_n869_), .A2(new_n240_), .A3(new_n472_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n856_), .A2(new_n473_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G183gat), .B1(new_n871_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1350gat));
  NAND2_X1  g678(.A1(new_n579_), .A2(new_n238_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n869_), .A2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n633_), .B(new_n857_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n882_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT125), .B1(new_n882_), .B2(G190gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n881_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT126), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n881_), .B(new_n887_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1351gat));
  NOR3_X1   g688(.A1(new_n376_), .A2(new_n649_), .A3(new_n383_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n803_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT127), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n803_), .A2(new_n893_), .A3(new_n890_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n436_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g696(.A(G204gat), .B1(new_n895_), .B2(new_n582_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n569_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n900_), .B2(new_n207_), .ZN(G1353gat));
  NAND2_X1  g700(.A1(new_n895_), .A2(new_n584_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT63), .B(G211gat), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n902_), .B2(new_n905_), .ZN(G1354gat));
  OAI21_X1  g705(.A(G218gat), .B1(new_n899_), .B2(new_n631_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n618_), .A2(G218gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n899_), .B2(new_n908_), .ZN(G1355gat));
endmodule


