//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT88), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT88), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n202_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT87), .Z(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT89), .ZN(new_n216_));
  INV_X1    g015(.A(new_n212_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT90), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n213_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n222_), .B(new_n223_), .C1(new_n217_), .C2(new_n218_), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n207_), .B(new_n210_), .C1(new_n220_), .C2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n216_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G127gat), .B(G134gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G113gat), .B(G120gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n227_), .B(new_n228_), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n229_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n216_), .A2(new_n231_), .A3(new_n225_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G225gat), .A2(G233gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(KEYINPUT100), .A3(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G1gat), .B(G29gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT0), .ZN(new_n237_));
  INV_X1    g036(.A(G57gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G85gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n230_), .A2(KEYINPUT4), .A3(new_n232_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n234_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n226_), .A2(new_n245_), .A3(new_n229_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n230_), .A2(new_n234_), .A3(new_n232_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT100), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n235_), .A2(new_n242_), .A3(new_n247_), .A4(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT33), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n242_), .B1(new_n233_), .B2(new_n244_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n243_), .A2(new_n234_), .A3(new_n246_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT101), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT101), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n258_), .A3(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n251_), .A2(new_n252_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n253_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT99), .ZN(new_n263_));
  INV_X1    g062(.A(G183gat), .ZN(new_n264_));
  INV_X1    g063(.A(G190gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT23), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT23), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(G183gat), .A3(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT79), .B(G190gat), .Z(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(G183gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT84), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT22), .ZN(new_n273_));
  OR3_X1    g072(.A1(new_n273_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n274_));
  INV_X1    g073(.A(G176gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(G169gat), .B1(new_n273_), .B2(KEYINPUT83), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT80), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n272_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n268_), .B(KEYINPUT82), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n266_), .A2(KEYINPUT81), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n266_), .A2(KEYINPUT81), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT25), .B(G183gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT26), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G190gat), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n285_), .B(new_n287_), .C1(new_n270_), .C2(new_n286_), .ZN(new_n288_));
  OR3_X1    g087(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n279_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n289_), .A3(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n284_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n280_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(G197gat), .B(G204gat), .Z(new_n297_));
  OAI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(KEYINPUT21), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT93), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n299_), .A3(KEYINPUT21), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n298_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n295_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT20), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT26), .B(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n285_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n291_), .A2(new_n278_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(new_n269_), .A4(new_n289_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n284_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT22), .B(G169gat), .Z(new_n309_));
  OAI21_X1  g108(.A(new_n279_), .B1(G176gat), .B2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n307_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n301_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n303_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n302_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT19), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(KEYINPUT98), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n311_), .A2(new_n312_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n316_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n280_), .A2(new_n294_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n312_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n319_), .A2(KEYINPUT20), .A3(new_n320_), .A4(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n320_), .B1(new_n302_), .B2(new_n313_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT98), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n318_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G64gat), .ZN(new_n330_));
  INV_X1    g129(.A(G92gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n263_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n332_), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT99), .B(new_n334_), .C1(new_n318_), .C2(new_n326_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n327_), .A2(new_n332_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n235_), .A2(new_n247_), .A3(new_n250_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n241_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n251_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n302_), .A2(new_n313_), .A3(new_n320_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT20), .B1(new_n311_), .B2(new_n312_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n343_), .B1(new_n312_), .B2(new_n321_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n342_), .B1(new_n344_), .B2(new_n320_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n318_), .A2(new_n326_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(new_n347_), .ZN(new_n350_));
  OAI22_X1  g149(.A1(new_n262_), .A2(new_n337_), .B1(new_n341_), .B2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n301_), .B1(new_n226_), .B2(KEYINPUT29), .ZN(new_n352_));
  AND2_X1   g151(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT94), .B(G233gat), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(G233gat), .B1(new_n353_), .B2(new_n354_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT94), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n352_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT96), .B1(new_n356_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n352_), .A2(new_n355_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT96), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n361_), .B(new_n362_), .C1(new_n352_), .C2(new_n358_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G78gat), .B(G106gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n364_), .B(KEYINPUT95), .Z(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT91), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT28), .B1(new_n226_), .B2(KEYINPUT29), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT28), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n216_), .A2(new_n369_), .A3(new_n370_), .A4(new_n225_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n367_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G22gat), .B(G50gat), .Z(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n374_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n375_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(new_n372_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n359_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n365_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n380_), .A2(new_n362_), .A3(new_n361_), .A4(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n366_), .A2(new_n376_), .A3(new_n379_), .A4(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n380_), .B(new_n361_), .C1(KEYINPUT97), .C2(new_n365_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n365_), .A2(KEYINPUT97), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n374_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n378_), .A2(new_n377_), .A3(new_n372_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n384_), .B(new_n386_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n321_), .B(KEYINPUT30), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n229_), .A2(KEYINPUT31), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n229_), .A2(KEYINPUT31), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n393_), .A2(KEYINPUT86), .A3(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n392_), .A2(KEYINPUT85), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n395_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n391_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n391_), .A2(new_n398_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G15gat), .B(G43gat), .Z(new_n402_));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n400_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n390_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n351_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT27), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n345_), .B2(new_n334_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n336_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n337_), .B2(new_n414_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n383_), .A2(new_n411_), .A3(new_n389_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n411_), .B1(new_n383_), .B2(new_n389_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n417_), .B(new_n341_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n413_), .A2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(G85gat), .A2(G92gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(G85gat), .A2(G92gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT66), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n240_), .A2(new_n331_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT66), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G85gat), .A2(G92gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n430_));
  NOR2_X1   g229(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n431_));
  OAI22_X1  g230(.A1(new_n430_), .A2(new_n431_), .B1(G99gat), .B2(G106gat), .ZN(new_n432_));
  AND3_X1   g231(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n436_));
  INV_X1    g235(.A(G99gat), .ZN(new_n437_));
  INV_X1    g236(.A(G106gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n429_), .A2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT64), .B1(new_n433_), .B2(new_n434_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G99gat), .A2(G106gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT64), .ZN(new_n446_));
  NAND3_X1  g245(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n442_), .A2(new_n448_), .A3(new_n432_), .A4(new_n439_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT8), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n424_), .A2(new_n428_), .A3(new_n450_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n441_), .A2(KEYINPUT8), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n442_), .A2(new_n448_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n425_), .A2(KEYINPUT9), .A3(new_n427_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(KEYINPUT9), .B2(new_n427_), .ZN(new_n455_));
  OR2_X1    g254(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n456_), .A2(new_n438_), .A3(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n453_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT67), .B1(new_n452_), .B2(new_n459_), .ZN(new_n460_));
  OR3_X1    g259(.A1(new_n453_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n451_), .A2(new_n449_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n450_), .B1(new_n429_), .B2(new_n440_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n461_), .B(new_n462_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G71gat), .B(G78gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(G57gat), .B(G64gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(KEYINPUT11), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  NAND3_X1  g269(.A1(new_n460_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n470_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n472_), .B(KEYINPUT12), .C1(new_n452_), .C2(new_n459_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n460_), .B2(new_n465_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n471_), .B(new_n473_), .C1(new_n474_), .C2(KEYINPUT12), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G230gat), .A2(G233gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n474_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n471_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n477_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G176gat), .B(G204gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(G120gat), .B(G148gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n478_), .A2(new_n481_), .A3(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n475_), .A2(new_n477_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n486_), .B(KEYINPUT69), .Z(new_n490_));
  OAI21_X1  g289(.A(new_n487_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT13), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n491_), .A2(KEYINPUT13), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G8gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT72), .B(G22gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G15gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT73), .B(G1gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT74), .B(G8gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n499_), .A2(G1gat), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G1gat), .ZN(new_n505_));
  INV_X1    g304(.A(G15gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n498_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n503_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n505_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n497_), .B1(new_n504_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(G1gat), .B1(new_n499_), .B2(new_n503_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(new_n508_), .A3(new_n505_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(G8gat), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G29gat), .B(G36gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G43gat), .B(G50gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT77), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n510_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n514_), .B2(new_n519_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n517_), .B(KEYINPUT15), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n510_), .A2(new_n526_), .A3(new_n513_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n522_), .A2(new_n524_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(G169gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(G197gat), .Z(new_n531_));
  OR2_X1    g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(KEYINPUT78), .A3(new_n531_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT78), .B1(new_n528_), .B2(new_n531_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n532_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n496_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n460_), .A2(new_n465_), .A3(new_n517_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n526_), .B1(new_n452_), .B2(new_n459_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT35), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G190gat), .B(G218gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(KEYINPUT36), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n538_), .A2(KEYINPUT71), .A3(new_n539_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT70), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n545_), .A2(new_n550_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n544_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n543_), .A2(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n544_), .A2(new_n551_), .A3(new_n556_), .A4(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT37), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n514_), .B(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(new_n470_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n470_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G127gat), .B(G155gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT76), .ZN(new_n567_));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT17), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n571_), .A2(KEYINPUT17), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n564_), .B(new_n565_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n565_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n572_), .B1(new_n576_), .B2(new_n563_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n558_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n560_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n537_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n421_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n340_), .B(KEYINPUT102), .Z(new_n585_));
  NOR3_X1   g384(.A1(new_n584_), .A2(new_n501_), .A3(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT38), .ZN(new_n587_));
  AOI211_X1 g386(.A(new_n340_), .B(new_n416_), .C1(new_n414_), .C2(new_n337_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n411_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n390_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n383_), .A2(new_n411_), .A3(new_n389_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n588_), .A2(new_n592_), .B1(new_n351_), .B2(new_n412_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n559_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n578_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n537_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n505_), .B1(new_n597_), .B2(new_n340_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n587_), .A2(new_n598_), .ZN(G1324gat));
  OR3_X1    g398(.A1(new_n584_), .A2(new_n417_), .A3(new_n502_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n417_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n594_), .A2(new_n601_), .A3(new_n596_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n602_), .A2(new_n603_), .A3(G8gat), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n602_), .B2(G8gat), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n600_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT103), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT103), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n600_), .B(new_n608_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n607_), .A2(KEYINPUT40), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT40), .B1(new_n607_), .B2(new_n609_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1325gat));
  AOI21_X1  g411(.A(new_n506_), .B1(new_n597_), .B2(new_n411_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT41), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n583_), .A2(new_n506_), .A3(new_n411_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1326gat));
  INV_X1    g415(.A(new_n390_), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n584_), .A2(G22gat), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n597_), .A2(new_n390_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(G22gat), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(KEYINPUT42), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(KEYINPUT42), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n618_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT104), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(KEYINPUT104), .B(new_n618_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1327gat));
  NOR2_X1   g426(.A1(new_n537_), .A2(new_n578_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n421_), .A2(new_n628_), .A3(new_n559_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n340_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n560_), .A2(new_n580_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n633_), .B2(KEYINPUT105), .ZN(new_n634_));
  INV_X1    g433(.A(new_n633_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n593_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n634_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n421_), .A2(new_n633_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(KEYINPUT44), .A3(new_n628_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n585_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(G29gat), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT44), .B1(new_n639_), .B2(new_n628_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n631_), .B1(new_n642_), .B2(new_n644_), .ZN(G1328gat));
  NAND2_X1  g444(.A1(new_n640_), .A2(new_n601_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G36gat), .B1(new_n646_), .B2(new_n643_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n629_), .A2(G36gat), .A3(new_n417_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT45), .Z(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1329gat));
  NAND3_X1  g451(.A1(new_n640_), .A2(G43gat), .A3(new_n411_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n629_), .A2(new_n589_), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n653_), .A2(new_n643_), .B1(G43gat), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g455(.A1(new_n640_), .A2(new_n390_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G50gat), .B1(new_n657_), .B2(new_n643_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n617_), .A2(G50gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT106), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n658_), .B1(new_n629_), .B2(new_n660_), .ZN(G1331gat));
  NOR3_X1   g460(.A1(new_n496_), .A2(new_n595_), .A3(new_n536_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n594_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n341_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n496_), .A2(new_n536_), .A3(new_n581_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n421_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n238_), .A3(new_n641_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(G1332gat));
  INV_X1    g468(.A(KEYINPUT48), .ZN(new_n670_));
  INV_X1    g469(.A(new_n663_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n601_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n672_), .B2(G64gat), .ZN(new_n673_));
  INV_X1    g472(.A(G64gat), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT48), .B(new_n674_), .C1(new_n671_), .C2(new_n601_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n601_), .A2(new_n674_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT107), .Z(new_n677_));
  OAI22_X1  g476(.A1(new_n673_), .A2(new_n675_), .B1(new_n666_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1333gat));
  OAI21_X1  g479(.A(G71gat), .B1(new_n663_), .B2(new_n589_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT49), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n589_), .A2(G71gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n666_), .B2(new_n683_), .ZN(G1334gat));
  OAI21_X1  g483(.A(G78gat), .B1(new_n663_), .B2(new_n617_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT50), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n617_), .A2(G78gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n666_), .B2(new_n687_), .ZN(G1335gat));
  NOR3_X1   g487(.A1(new_n496_), .A2(new_n578_), .A3(new_n536_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n593_), .A2(new_n690_), .A3(new_n558_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n240_), .A3(new_n641_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n593_), .A2(new_n635_), .A3(new_n634_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n637_), .B1(new_n421_), .B2(new_n633_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n689_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT109), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n639_), .A2(new_n697_), .A3(new_n689_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n341_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n692_), .B1(new_n699_), .B2(new_n240_), .ZN(G1336gat));
  AOI21_X1  g499(.A(G92gat), .B1(new_n691_), .B2(new_n601_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT110), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n696_), .A2(new_n698_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n417_), .A2(new_n331_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(G1337gat));
  OR2_X1    g504(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n706_));
  NAND2_X1  g505(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n437_), .B1(new_n703_), .B2(new_n411_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n691_), .A2(new_n456_), .A3(new_n457_), .A4(new_n411_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n706_), .B(new_n707_), .C1(new_n708_), .C2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n697_), .B1(new_n639_), .B2(new_n689_), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT109), .B(new_n690_), .C1(new_n636_), .C2(new_n638_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n411_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G99gat), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n715_), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n709_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n711_), .A2(new_n716_), .ZN(G1338gat));
  OAI211_X1 g516(.A(new_n390_), .B(new_n689_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n639_), .A2(KEYINPUT112), .A3(new_n390_), .A4(new_n689_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n438_), .B1(new_n722_), .B2(KEYINPUT52), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(KEYINPUT52), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n725_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .A4(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n691_), .A2(new_n438_), .A3(new_n390_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT53), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT53), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n726_), .A2(new_n732_), .A3(new_n728_), .A4(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1339gat));
  NOR2_X1   g533(.A1(new_n585_), .A2(new_n601_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n418_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT57), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n522_), .A2(new_n523_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n531_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n520_), .A2(new_n524_), .A3(new_n527_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n522_), .A2(new_n524_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n525_), .A2(new_n527_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n531_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT78), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n742_), .B1(new_n747_), .B2(new_n533_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n491_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT114), .B1(new_n475_), .B2(new_n477_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT55), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT114), .B(new_n752_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n475_), .A2(new_n477_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n490_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(KEYINPUT56), .A3(new_n756_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n750_), .A2(KEYINPUT55), .B1(new_n477_), .B2(new_n475_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n490_), .B1(new_n758_), .B2(new_n753_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n536_), .A2(new_n487_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n749_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n737_), .B1(new_n763_), .B2(new_n559_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n747_), .A2(new_n533_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n765_), .A2(new_n487_), .A3(new_n741_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n767_), .B(new_n490_), .C1(new_n758_), .C2(new_n753_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n755_), .B2(new_n756_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT58), .B(new_n766_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n633_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n536_), .A2(new_n487_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n755_), .A2(new_n756_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n760_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n775_), .B1(new_n778_), .B2(new_n757_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT57), .B(new_n558_), .C1(new_n779_), .C2(new_n749_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n764_), .A2(new_n774_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n595_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n494_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n536_), .B1(new_n783_), .B2(new_n492_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT54), .B1(new_n785_), .B2(new_n581_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n635_), .A2(new_n784_), .A3(new_n787_), .A4(new_n578_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n736_), .B1(new_n782_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G113gat), .B1(new_n790_), .B2(new_n536_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT116), .Z(new_n792_));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n790_), .B2(new_n794_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n781_), .A2(new_n595_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT117), .B(KEYINPUT59), .C1(new_n796_), .C2(new_n736_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n790_), .B2(new_n794_), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n796_), .A2(KEYINPUT118), .A3(KEYINPUT59), .A4(new_n736_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT119), .B1(new_n798_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n790_), .A2(new_n794_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT118), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n790_), .A2(new_n799_), .A3(new_n794_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n795_), .A2(new_n797_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n803_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n536_), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT120), .B(G113gat), .Z(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n792_), .B1(new_n811_), .B2(new_n814_), .ZN(G1340gat));
  INV_X1    g614(.A(G120gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n496_), .B2(KEYINPUT60), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n790_), .B(new_n817_), .C1(KEYINPUT60), .C2(new_n816_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT121), .Z(new_n819_));
  NOR3_X1   g618(.A1(new_n798_), .A2(new_n802_), .A3(new_n496_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n816_), .ZN(G1341gat));
  AOI21_X1  g620(.A(G127gat), .B1(new_n790_), .B2(new_n578_), .ZN(new_n822_));
  INV_X1    g621(.A(G127gat), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(KEYINPUT122), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n578_), .A2(G127gat), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(KEYINPUT122), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n822_), .B1(new_n811_), .B2(new_n826_), .ZN(G1342gat));
  INV_X1    g626(.A(G134gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n790_), .A2(new_n828_), .A3(new_n559_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n635_), .B1(new_n803_), .B2(new_n810_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n828_), .ZN(G1343gat));
  NOR4_X1   g630(.A1(new_n796_), .A2(new_n590_), .A3(new_n601_), .A4(new_n585_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n536_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n495_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g635(.A1(new_n796_), .A2(new_n590_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n578_), .A3(new_n735_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(KEYINPUT123), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n832_), .B2(new_n578_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT61), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n838_), .A2(KEYINPUT123), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n832_), .A2(new_n840_), .A3(new_n578_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT61), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n842_), .A2(G155gat), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G155gat), .B1(new_n842_), .B2(new_n846_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1346gat));
  INV_X1    g648(.A(new_n832_), .ZN(new_n850_));
  OR3_X1    g649(.A1(new_n850_), .A2(G162gat), .A3(new_n558_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G162gat), .B1(new_n850_), .B2(new_n635_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1347gat));
  NOR2_X1   g652(.A1(new_n796_), .A2(new_n390_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n641_), .A2(new_n589_), .A3(new_n417_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n536_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(G169gat), .A3(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n309_), .B2(new_n858_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n858_), .B2(G169gat), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1348gat));
  AOI21_X1  g662(.A(G176gat), .B1(new_n857_), .B2(new_n495_), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n854_), .B(KEYINPUT125), .Z(new_n865_));
  AND3_X1   g664(.A1(new_n855_), .A2(G176gat), .A3(new_n495_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  NOR3_X1   g666(.A1(new_n856_), .A2(new_n285_), .A3(new_n595_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n578_), .A3(new_n855_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n264_), .ZN(G1350gat));
  OAI21_X1  g669(.A(G190gat), .B1(new_n856_), .B2(new_n635_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n559_), .A2(new_n304_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n856_), .B2(new_n872_), .ZN(G1351gat));
  NOR2_X1   g672(.A1(new_n417_), .A2(new_n340_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n837_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n812_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT126), .B(G197gat), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1352gat));
  INV_X1    g677(.A(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n495_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n578_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n883_));
  AND2_X1   g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n882_), .B2(new_n883_), .ZN(G1354gat));
  AOI21_X1  g685(.A(G218gat), .B1(new_n879_), .B2(new_n559_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n633_), .A2(G218gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT127), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n879_), .B2(new_n889_), .ZN(G1355gat));
endmodule


