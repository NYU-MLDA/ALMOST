//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT86), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n209_), .A3(KEYINPUT1), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G155gat), .ZN(new_n212_));
  INV_X1    g011(.A(G162gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT85), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(G155gat), .B2(G162gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G155gat), .A3(G162gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n205_), .B1(new_n211_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(new_n216_), .A3(new_n206_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  INV_X1    g023(.A(G141gat), .ZN(new_n225_));
  INV_X1    g024(.A(G148gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n202_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n227_), .A2(new_n229_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n223_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n220_), .A2(new_n221_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT87), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT87), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n220_), .A2(new_n233_), .A3(new_n236_), .A4(new_n221_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G22gat), .B(G50gat), .Z(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n235_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n242_));
  XOR2_X1   g041(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n235_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n239_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n243_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G228gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n221_), .B1(new_n220_), .B2(new_n233_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT21), .ZN(new_n252_));
  INV_X1    g051(.A(G218gat), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n253_), .A2(G211gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(G211gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n252_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT21), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n259_), .A3(KEYINPUT21), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n250_), .B1(new_n251_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n205_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n206_), .A2(new_n209_), .A3(KEYINPUT1), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n209_), .B1(new_n206_), .B2(KEYINPUT1), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n214_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n266_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n227_), .A2(new_n231_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n229_), .A2(new_n230_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n222_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT29), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(new_n249_), .A3(new_n263_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G78gat), .B(G106gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n265_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT91), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT91), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n265_), .A2(new_n276_), .A3(new_n281_), .A4(new_n278_), .ZN(new_n282_));
  AND4_X1   g081(.A1(new_n245_), .A2(new_n248_), .A3(new_n280_), .A4(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n265_), .A2(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n277_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT90), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n248_), .A2(new_n245_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n279_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(KEYINPUT89), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT89), .B1(new_n289_), .B2(new_n290_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n288_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT83), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G169gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT22), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT22), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT22), .B(G169gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT81), .A3(new_n309_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n304_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n318_), .B2(new_n303_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT25), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n323_));
  INV_X1    g122(.A(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT26), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G190gat), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n321_), .A2(new_n323_), .A3(new_n325_), .A4(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n319_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT82), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n315_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n312_), .A2(new_n314_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n331_), .A2(new_n300_), .B1(G169gat), .B2(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n319_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT82), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n296_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341_));
  INV_X1    g140(.A(G43gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G15gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n343_), .B(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n333_), .B1(new_n315_), .B2(new_n332_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n337_), .A2(KEYINPUT82), .A3(new_n338_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT30), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n340_), .A2(new_n346_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n346_), .B1(new_n340_), .B2(new_n349_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n295_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n346_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n349_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT30), .B1(new_n347_), .B2(new_n348_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n340_), .A2(new_n346_), .A3(new_n349_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(KEYINPUT83), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G134gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G127gat), .ZN(new_n360_));
  INV_X1    g159(.A(G113gat), .ZN(new_n361_));
  INV_X1    g160(.A(G120gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(G127gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G134gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G113gat), .A2(G120gat), .ZN(new_n366_));
  AND4_X1   g165(.A1(new_n360_), .A2(new_n363_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n360_), .A2(new_n365_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT31), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n352_), .A2(new_n358_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n295_), .B(new_n372_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT84), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n376_), .A3(new_n373_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n294_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n347_), .A2(new_n348_), .A3(new_n264_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n336_), .A2(new_n310_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n325_), .A2(new_n327_), .ZN(new_n382_));
  XOR2_X1   g181(.A(KEYINPUT25), .B(G183gat), .Z(new_n383_));
  OAI211_X1 g182(.A(new_n319_), .B(new_n331_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n380_), .B1(new_n385_), .B2(new_n263_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT19), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT20), .B1(new_n385_), .B2(new_n263_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n389_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n334_), .A2(new_n339_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(new_n393_), .C1(new_n394_), .C2(new_n264_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(G64gat), .B(G92gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n396_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n396_), .A2(new_n402_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n367_), .A2(new_n368_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n220_), .A2(new_n233_), .A3(new_n369_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n369_), .B1(new_n220_), .B2(new_n233_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n407_), .A2(KEYINPUT4), .A3(new_n408_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT93), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT93), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n411_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT0), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G57gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G85gat), .ZN(new_n425_));
  INV_X1    g224(.A(G57gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n423_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G85gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n420_), .A2(KEYINPUT33), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n430_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n415_), .B(new_n409_), .C1(KEYINPUT4), .C2(new_n407_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n407_), .A2(new_n408_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n432_), .B(new_n433_), .C1(new_n434_), .C2(new_n409_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n404_), .A2(new_n405_), .A3(new_n431_), .A4(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT94), .B1(new_n420_), .B2(new_n430_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n414_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n418_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n410_), .B(new_n430_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT94), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n437_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT95), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n420_), .A2(KEYINPUT94), .A3(new_n430_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(new_n442_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(KEYINPUT95), .A3(new_n437_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n436_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n420_), .A2(new_n430_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n441_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n392_), .B1(new_n394_), .B2(new_n264_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n389_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT96), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n379_), .A2(KEYINPUT96), .A3(new_n393_), .A4(new_n386_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(KEYINPUT32), .A3(new_n401_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n390_), .A2(new_n395_), .A3(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n453_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n378_), .B1(new_n451_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n453_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467_));
  INV_X1    g266(.A(new_n405_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n468_), .B2(new_n403_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n459_), .A2(new_n402_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n404_), .A2(new_n470_), .A3(KEYINPUT27), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n246_), .A2(new_n247_), .A3(new_n243_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n244_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n290_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n478_), .A2(new_n291_), .B1(new_n287_), .B2(new_n283_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n294_), .A2(new_n374_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n473_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n465_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT67), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G120gat), .B(G148gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT5), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G176gat), .B(G204gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G71gat), .B(G78gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT11), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n492_));
  INV_X1    g291(.A(new_n490_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n491_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G85gat), .B(G92gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT9), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT10), .B(G99gat), .Z(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(G85gat), .A3(G92gat), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n499_), .A2(new_n502_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n497_), .A2(KEYINPUT64), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511_));
  INV_X1    g310(.A(G99gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n501_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n513_), .A2(new_n505_), .A3(new_n506_), .A4(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n510_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n510_), .B2(new_n515_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n496_), .B(new_n509_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT12), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n509_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n496_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT65), .B1(new_n518_), .B2(new_n519_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n519_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT65), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n517_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n529_), .A3(new_n509_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n523_), .A2(KEYINPUT12), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n525_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n524_), .A2(new_n520_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(G230gat), .A3(G233gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n536_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n484_), .B(new_n488_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n488_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(new_n539_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n535_), .A2(new_n538_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT67), .B1(new_n547_), .B2(new_n543_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n542_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT13), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n542_), .B(KEYINPUT13), .C1(new_n545_), .C2(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(G1gat), .ZN(new_n554_));
  INV_X1    g353(.A(G8gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G22gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(G15gat), .ZN(new_n558_));
  INV_X1    g357(.A(G15gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(G22gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT74), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G1gat), .B(G8gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n561_), .A2(KEYINPUT74), .ZN(new_n565_));
  INV_X1    g364(.A(new_n563_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(KEYINPUT74), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G36gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(G29gat), .ZN(new_n571_));
  INV_X1    g370(.A(G29gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(G36gat), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n571_), .A2(new_n573_), .A3(KEYINPUT69), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT69), .B1(new_n571_), .B2(new_n573_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT70), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n573_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT70), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n571_), .A2(new_n573_), .A3(KEYINPUT69), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G43gat), .B(G50gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n576_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n583_), .B1(new_n576_), .B2(new_n582_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n569_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n576_), .A2(new_n582_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n583_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n564_), .A2(new_n590_), .A3(new_n584_), .A4(new_n568_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT77), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(KEYINPUT77), .A3(new_n591_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n585_), .A2(new_n586_), .A3(KEYINPUT15), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT15), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n590_), .B2(new_n584_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n568_), .B(new_n564_), .C1(new_n599_), .C2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n587_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n595_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G169gat), .B(G197gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT79), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT79), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n598_), .A2(new_n604_), .A3(new_n610_), .A4(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n598_), .A2(new_n604_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n607_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT78), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n612_), .A2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n609_), .A2(new_n615_), .A3(new_n616_), .A4(new_n611_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n553_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n483_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT35), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n522_), .B1(new_n584_), .B2(new_n590_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT15), .B1(new_n585_), .B2(new_n586_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n590_), .A2(new_n600_), .A3(new_n584_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n631_), .B2(new_n530_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n627_), .B1(new_n632_), .B2(KEYINPUT71), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n530_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n628_), .ZN(new_n635_));
  AND4_X1   g434(.A1(KEYINPUT71), .A2(new_n634_), .A3(new_n635_), .A4(new_n627_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n624_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n635_), .A3(KEYINPUT71), .ZN(new_n638_));
  INV_X1    g437(.A(new_n627_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n632_), .A2(KEYINPUT71), .A3(new_n627_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n632_), .A2(new_n624_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(G190gat), .B(G218gat), .Z(new_n644_));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT36), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n637_), .A2(new_n643_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT72), .B1(new_n637_), .B2(new_n643_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n647_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n651_), .ZN(new_n653_));
  AOI211_X1 g452(.A(KEYINPUT72), .B(new_n653_), .C1(new_n637_), .C2(new_n643_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n623_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT72), .ZN(new_n656_));
  INV_X1    g455(.A(new_n643_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT35), .B1(new_n640_), .B2(new_n641_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n656_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n653_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n650_), .A2(new_n651_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT73), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(KEYINPUT37), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n649_), .A4(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n655_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(G231gat), .A2(G233gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n496_), .B(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(new_n569_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(G127gat), .B(G155gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(G183gat), .B(G211gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT17), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n668_), .A2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n673_), .B(KEYINPUT17), .Z(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(new_n668_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT76), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n665_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n622_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n554_), .A3(new_n453_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT97), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT38), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT99), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n652_), .A2(new_n654_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n465_), .B2(new_n482_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n678_), .A3(new_n621_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G1gat), .B1(new_n690_), .B2(new_n466_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n683_), .A2(new_n684_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(KEYINPUT98), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT98), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n683_), .A2(new_n694_), .A3(new_n684_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n686_), .B(new_n691_), .C1(new_n693_), .C2(new_n695_), .ZN(G1324gat));
  NAND2_X1  g495(.A1(new_n471_), .A2(new_n469_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G8gat), .B1(new_n690_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT39), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n681_), .A2(new_n555_), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(G1325gat));
  INV_X1    g503(.A(new_n377_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n376_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G15gat), .B1(new_n690_), .B2(new_n708_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(KEYINPUT41), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(KEYINPUT41), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n681_), .A2(new_n559_), .A3(new_n707_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(G1326gat));
  OAI21_X1  g512(.A(G22gat), .B1(new_n690_), .B2(new_n479_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n715_));
  OR2_X1    g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n715_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n681_), .A2(new_n557_), .A3(new_n294_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n716_), .A2(new_n717_), .A3(new_n718_), .ZN(G1327gat));
  NOR2_X1   g518(.A1(new_n687_), .A2(new_n678_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n622_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT104), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n622_), .A2(new_n723_), .A3(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G29gat), .B1(new_n726_), .B2(new_n453_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n553_), .A2(new_n620_), .A3(new_n678_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n483_), .A2(new_n730_), .A3(new_n665_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n483_), .B2(new_n665_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n728_), .B(new_n729_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT44), .B1(new_n733_), .B2(KEYINPUT103), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT102), .B1(KEYINPUT103), .B2(KEYINPUT44), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n483_), .A2(new_n665_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT43), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n483_), .A2(new_n665_), .A3(new_n730_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n735_), .B1(new_n739_), .B2(new_n729_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n734_), .A2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n466_), .A2(new_n572_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n727_), .B1(new_n741_), .B2(new_n742_), .ZN(G1328gat));
  NAND2_X1  g542(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n697_), .B1(new_n734_), .B2(new_n740_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G36gat), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT105), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n748_), .A3(G36gat), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n697_), .B(KEYINPUT106), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n722_), .A2(new_n570_), .A3(new_n724_), .A4(new_n753_), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n755_));
  OR2_X1    g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n755_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n751_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n744_), .B1(new_n750_), .B2(new_n758_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n745_), .A2(new_n748_), .A3(G36gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n748_), .B1(new_n745_), .B2(G36gat), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n758_), .B(new_n744_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n759_), .A2(new_n763_), .ZN(G1329gat));
  NOR3_X1   g563(.A1(new_n725_), .A2(G43gat), .A3(new_n708_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n374_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n741_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n767_), .B2(G43gat), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g568(.A1(new_n741_), .A2(new_n294_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n770_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT109), .B1(new_n770_), .B2(G50gat), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n479_), .A2(G50gat), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT110), .Z(new_n774_));
  OAI22_X1  g573(.A1(new_n771_), .A2(new_n772_), .B1(new_n725_), .B2(new_n774_), .ZN(G1331gat));
  INV_X1    g574(.A(new_n553_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n620_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(new_n483_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(new_n680_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n426_), .A3(new_n453_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n689_), .A2(new_n778_), .A3(new_n678_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G57gat), .B1(new_n782_), .B2(new_n466_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1332gat));
  OAI21_X1  g583(.A(G64gat), .B1(new_n782_), .B2(new_n752_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT48), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n752_), .A2(G64gat), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT111), .Z(new_n788_));
  NAND2_X1  g587(.A1(new_n780_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(G1333gat));
  OAI21_X1  g589(.A(G71gat), .B1(new_n782_), .B2(new_n708_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT49), .ZN(new_n792_));
  INV_X1    g591(.A(G71gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n780_), .A2(new_n793_), .A3(new_n707_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1334gat));
  OAI21_X1  g594(.A(G78gat), .B1(new_n782_), .B2(new_n479_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT50), .ZN(new_n797_));
  INV_X1    g596(.A(G78gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n780_), .A2(new_n798_), .A3(new_n294_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1335gat));
  NAND2_X1  g599(.A1(new_n779_), .A2(new_n720_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(new_n428_), .A3(new_n453_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n776_), .A2(new_n678_), .A3(new_n777_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n739_), .A2(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n805_), .A2(new_n453_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n803_), .B1(new_n806_), .B2(new_n428_), .ZN(G1336gat));
  INV_X1    g606(.A(G92gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n802_), .A2(new_n808_), .A3(new_n697_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n805_), .A2(new_n753_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n808_), .ZN(G1337gat));
  AOI21_X1  g610(.A(new_n512_), .B1(new_n805_), .B2(new_n707_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n766_), .A2(new_n500_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n802_), .B2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(G1338gat));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n739_), .A2(new_n294_), .A3(new_n804_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G106gat), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(KEYINPUT113), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(KEYINPUT113), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n817_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n819_), .A2(KEYINPUT113), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(KEYINPUT113), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(KEYINPUT52), .A3(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n802_), .A2(new_n501_), .A3(new_n294_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n822_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g627(.A1(new_n777_), .A2(new_n553_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(new_n655_), .A3(new_n664_), .A4(new_n678_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n547_), .A2(new_n543_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n603_), .A2(KEYINPUT115), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n602_), .B2(new_n587_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n596_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n594_), .A2(new_n597_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n614_), .B1(new_n839_), .B2(new_n595_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n838_), .A2(new_n840_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n525_), .A2(new_n533_), .A3(KEYINPUT55), .A4(new_n534_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT114), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n530_), .A2(new_n532_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(KEYINPUT55), .A4(new_n534_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n534_), .B1(new_n525_), .B2(new_n533_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n535_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n543_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(KEYINPUT56), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n853_), .B(new_n543_), .C1(new_n847_), .C2(new_n850_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n834_), .B(new_n841_), .C1(new_n852_), .C2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT118), .B1(new_n855_), .B2(KEYINPUT117), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n857_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n856_), .A2(new_n857_), .B1(new_n855_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n665_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n833_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n851_), .B(KEYINPUT56), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n864_), .A2(new_n858_), .A3(new_n834_), .A4(new_n841_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT58), .B1(new_n865_), .B2(KEYINPUT118), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n855_), .A2(new_n860_), .ZN(new_n867_));
  OAI211_X1 g666(.A(KEYINPUT119), .B(new_n665_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n549_), .A2(new_n841_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n549_), .A2(KEYINPUT116), .A3(new_n841_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n834_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n620_), .A2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(KEYINPUT57), .B(new_n687_), .C1(new_n873_), .C2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n687_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n863_), .A2(new_n868_), .A3(new_n876_), .A4(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n832_), .B1(new_n880_), .B2(new_n679_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n698_), .A2(new_n479_), .A3(new_n766_), .A4(new_n453_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT120), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT121), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n679_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n832_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n883_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n885_), .A2(new_n890_), .A3(new_n777_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n361_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(new_n361_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n888_), .B2(new_n883_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n884_), .A2(KEYINPUT59), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n665_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n879_), .A3(KEYINPUT123), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n876_), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT123), .B1(new_n899_), .B2(new_n879_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n679_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n898_), .B1(new_n903_), .B2(new_n887_), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n896_), .A2(new_n904_), .A3(new_n361_), .A4(new_n620_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n893_), .A2(new_n894_), .A3(new_n905_), .ZN(G1340gat));
  NOR2_X1   g705(.A1(new_n896_), .A2(new_n904_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G120gat), .B1(new_n908_), .B2(new_n776_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n885_), .A2(new_n890_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n553_), .A2(new_n911_), .A3(new_n362_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n911_), .B2(new_n362_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n909_), .A2(new_n914_), .ZN(G1341gat));
  OAI21_X1  g714(.A(G127gat), .B1(new_n908_), .B2(new_n679_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n910_), .A2(new_n364_), .A3(new_n678_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1342gat));
  AOI21_X1  g717(.A(G134gat), .B1(new_n910_), .B2(new_n688_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n665_), .A2(G134gat), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(KEYINPUT124), .Z(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n907_), .B2(new_n921_), .ZN(G1343gat));
  OAI21_X1  g721(.A(new_n294_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n881_), .A2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n924_), .A2(new_n453_), .A3(new_n752_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n620_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n225_), .ZN(G1344gat));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n776_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT125), .B(G148gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1345gat));
  NOR2_X1   g729(.A1(new_n925_), .A2(new_n679_), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT61), .B(G155gat), .Z(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1346gat));
  OAI21_X1  g732(.A(G162gat), .B1(new_n925_), .B2(new_n862_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n688_), .A2(new_n213_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n925_), .B2(new_n935_), .ZN(G1347gat));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n903_), .A2(new_n887_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n752_), .A2(new_n453_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n707_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n294_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n620_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n937_), .B1(new_n943_), .B2(new_n305_), .ZN(new_n944_));
  OAI211_X1 g743(.A(KEYINPUT62), .B(G169gat), .C1(new_n942_), .C2(new_n620_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n313_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n944_), .A2(new_n945_), .A3(new_n946_), .ZN(G1348gat));
  NAND3_X1  g746(.A1(new_n938_), .A2(new_n553_), .A3(new_n941_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n881_), .A2(new_n294_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n940_), .A2(new_n309_), .A3(new_n776_), .ZN(new_n950_));
  AOI22_X1  g749(.A1(new_n948_), .A2(new_n309_), .B1(new_n949_), .B2(new_n950_), .ZN(G1349gat));
  NAND4_X1  g750(.A1(new_n938_), .A2(new_n678_), .A3(new_n383_), .A4(new_n941_), .ZN(new_n952_));
  NOR4_X1   g751(.A1(new_n881_), .A2(new_n679_), .A3(new_n294_), .A4(new_n940_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n953_), .B2(G183gat), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  OAI211_X1 g755(.A(new_n952_), .B(KEYINPUT126), .C1(new_n953_), .C2(G183gat), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1350gat));
  OAI21_X1  g757(.A(G190gat), .B1(new_n942_), .B2(new_n862_), .ZN(new_n959_));
  OR2_X1    g758(.A1(new_n687_), .A2(new_n382_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n942_), .B2(new_n960_), .ZN(G1351gat));
  AND2_X1   g760(.A1(new_n924_), .A2(new_n939_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(new_n777_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g763(.A1(new_n962_), .A2(KEYINPUT127), .A3(G204gat), .A4(new_n553_), .ZN(new_n965_));
  XOR2_X1   g764(.A(KEYINPUT127), .B(G204gat), .Z(new_n966_));
  NAND2_X1  g765(.A1(new_n924_), .A2(new_n939_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n967_), .B2(new_n776_), .ZN(new_n968_));
  AND2_X1   g767(.A1(new_n965_), .A2(new_n968_), .ZN(G1353gat));
  AOI21_X1  g768(.A(new_n679_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n970_));
  AND3_X1   g769(.A1(new_n924_), .A2(new_n939_), .A3(new_n970_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1354gat));
  NAND3_X1  g772(.A1(new_n962_), .A2(new_n253_), .A3(new_n688_), .ZN(new_n974_));
  OAI21_X1  g773(.A(G218gat), .B1(new_n967_), .B2(new_n862_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n974_), .A2(new_n975_), .ZN(G1355gat));
endmodule


