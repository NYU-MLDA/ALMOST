//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT25), .B(G183gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT80), .B(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT26), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n212_), .B1(G169gat), .B2(G176gat), .ZN(new_n213_));
  NOR3_X1   g012(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n216_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n220_));
  OAI22_X1  g019(.A1(new_n218_), .A2(KEYINPUT23), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n211_), .A2(new_n215_), .A3(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(KEYINPUT23), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT83), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n219_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n218_), .A2(new_n229_), .A3(KEYINPUT23), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G183gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n207_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n225_), .B1(new_n234_), .B2(KEYINPUT84), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT84), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n231_), .A2(new_n236_), .A3(new_n233_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n222_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G204gat), .ZN(new_n240_));
  INV_X1    g039(.A(G204gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G197gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT21), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT95), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G211gat), .B(G218gat), .Z(new_n247_));
  INV_X1    g046(.A(KEYINPUT94), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n240_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n239_), .A2(KEYINPUT94), .A3(G204gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n242_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n247_), .B1(new_n251_), .B2(KEYINPUT21), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n247_), .A2(KEYINPUT21), .A3(new_n243_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT20), .B1(new_n238_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n206_), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT26), .B(G190gat), .Z(new_n259_));
  OAI211_X1 g058(.A(new_n231_), .B(new_n215_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n221_), .B1(G183gat), .B2(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n224_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(new_n255_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n205_), .B1(new_n257_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n238_), .A2(new_n256_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n263_), .B2(new_n255_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n204_), .A3(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT18), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  AOI22_X1  g072(.A1(new_n265_), .A2(new_n269_), .B1(KEYINPUT32), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT98), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n263_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n260_), .A2(KEYINPUT98), .A3(new_n262_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n256_), .A3(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n278_), .B(KEYINPUT20), .C1(new_n256_), .C2(new_n238_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n204_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n266_), .A2(new_n268_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n205_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n273_), .A2(KEYINPUT32), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n274_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G1gat), .B(G29gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(G85gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT0), .B(G57gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT86), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT1), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n295_), .B2(KEYINPUT1), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n296_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n299_), .B2(new_n298_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n304_), .B(KEYINPUT2), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n302_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT3), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT89), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n309_), .A2(new_n314_), .A3(KEYINPUT89), .A4(new_n312_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n295_), .B1(G155gat), .B2(G162gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT90), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n323_));
  AOI211_X1 g122(.A(new_n323_), .B(new_n320_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n305_), .B(new_n308_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n305_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n308_), .B(KEYINPUT85), .ZN(new_n328_));
  OAI211_X1 g127(.A(KEYINPUT4), .B(new_n325_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330_));
  INV_X1    g129(.A(new_n328_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n326_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT97), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n325_), .B(new_n333_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n290_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n336_), .A3(new_n290_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT99), .A3(new_n339_), .ZN(new_n340_));
  AOI211_X1 g139(.A(KEYINPUT99), .B(new_n290_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n286_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n273_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n265_), .A2(new_n269_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT33), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n339_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n329_), .A2(new_n333_), .A3(new_n332_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n290_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n325_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n334_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n350_), .B(new_n351_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n339_), .A2(new_n348_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n347_), .A2(new_n349_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n343_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G78gat), .B(G106gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n326_), .A2(KEYINPUT29), .ZN(new_n359_));
  INV_X1    g158(.A(G228gat), .ZN(new_n360_));
  INV_X1    g159(.A(G233gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n256_), .A2(KEYINPUT93), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n359_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n359_), .B2(new_n364_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n358_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT96), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n322_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n324_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n372_), .A2(new_n373_), .A3(new_n305_), .A4(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n374_), .B1(new_n326_), .B2(KEYINPUT29), .ZN(new_n377_));
  XOR2_X1   g176(.A(G22gat), .B(G50gat), .Z(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n359_), .A2(new_n364_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n362_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n359_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n358_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(KEYINPUT96), .B(new_n358_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n369_), .A2(new_n382_), .A3(new_n387_), .A4(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n367_), .A2(new_n387_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n381_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(KEYINPUT92), .A3(new_n379_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(G15gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT30), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n238_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n238_), .A2(new_n400_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n328_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405_));
  INV_X1    g204(.A(G43gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT31), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n238_), .A2(new_n400_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(new_n331_), .A3(new_n401_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n404_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n404_), .B2(new_n410_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n396_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n357_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n346_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n283_), .A2(new_n344_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n416_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n339_), .A2(KEYINPUT99), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n422_), .A2(new_n337_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT100), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n341_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT100), .B1(new_n340_), .B2(new_n342_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n421_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n411_), .A2(new_n412_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n396_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n413_), .A2(new_n389_), .A3(new_n395_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n415_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(G85gat), .A2(G92gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G85gat), .A2(G92gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G99gat), .A2(G106gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT6), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(G99gat), .A3(G106gat), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n435_), .A2(KEYINPUT9), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n441_));
  INV_X1    g240(.A(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT9), .ZN(new_n445_));
  INV_X1    g244(.A(G85gat), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n446_), .A2(KEYINPUT64), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(KEYINPUT64), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n445_), .B(G92gat), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n440_), .A2(KEYINPUT65), .A3(new_n444_), .A4(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT65), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT64), .B(G85gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n445_), .A2(G92gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n444_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n437_), .A2(new_n439_), .ZN(new_n455_));
  INV_X1    g254(.A(G92gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n446_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(KEYINPUT9), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n451_), .B1(new_n454_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n435_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT7), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G99gat), .A2(G106gat), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n437_), .A2(new_n439_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT66), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT66), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n468_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n462_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT8), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI211_X1 g272(.A(KEYINPUT8), .B(new_n462_), .C1(new_n465_), .C2(new_n470_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n450_), .B(new_n461_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(G29gat), .B(G36gat), .Z(new_n477_));
  XOR2_X1   g276(.A(G43gat), .B(G50gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G232gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n476_), .A2(new_n479_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n467_), .A2(new_n469_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n464_), .A2(new_n463_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n438_), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n436_), .A2(KEYINPUT6), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n435_), .B1(new_n485_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT8), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n471_), .A2(new_n472_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n461_), .A2(new_n450_), .A3(KEYINPUT69), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT69), .B1(new_n461_), .B2(new_n450_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n479_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT15), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n479_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n484_), .A2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n483_), .A2(new_n480_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(KEYINPUT36), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n507_), .B(KEYINPUT36), .Z(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n504_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n432_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G64gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G57gat), .ZN(new_n518_));
  INV_X1    g317(.A(G57gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(G64gat), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT11), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G71gat), .B(G78gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT67), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G71gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G78gat), .ZN(new_n525_));
  INV_X1    g324(.A(G78gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G71gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n528_), .B(new_n529_), .C1(new_n530_), .C2(KEYINPUT11), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(KEYINPUT11), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n523_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n523_), .B2(new_n531_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT11), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n519_), .A2(G64gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n517_), .A2(G57gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n529_), .B1(new_n541_), .B2(new_n528_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n521_), .A2(KEYINPUT67), .A3(new_n522_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n532_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n523_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT68), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n537_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n534_), .A2(new_n535_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n547_), .A2(new_n476_), .B1(new_n496_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n536_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n544_), .A2(KEYINPUT68), .A3(new_n545_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n461_), .A2(new_n450_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n553_), .A2(new_n554_), .B1(new_n493_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n552_), .B1(new_n556_), .B2(KEYINPUT12), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n475_), .B1(new_n537_), .B2(new_n546_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT70), .A3(new_n549_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n551_), .A2(new_n557_), .A3(new_n559_), .A4(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n475_), .A2(new_n537_), .A3(new_n546_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n563_), .B2(new_n556_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G120gat), .B(G148gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n561_), .A2(new_n564_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT72), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(KEYINPUT72), .A3(new_n573_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(KEYINPUT13), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n571_), .A2(KEYINPUT72), .A3(new_n573_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n579_), .B2(new_n574_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT74), .B(G8gat), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT14), .B1(new_n581_), .B2(new_n202_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G15gat), .B(G22gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G1gat), .B(G8gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n583_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n498_), .A2(new_n585_), .A3(new_n588_), .A4(new_n500_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n479_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n589_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n590_), .B(new_n497_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n593_), .B1(new_n594_), .B2(new_n592_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT79), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G113gat), .B(G141gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(G169gat), .B(G197gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n597_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n595_), .A2(new_n596_), .A3(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n607_));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n590_), .B(new_n612_), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n548_), .B(KEYINPUT75), .ZN(new_n615_));
  AOI211_X1 g414(.A(new_n607_), .B(new_n611_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n611_), .B(KEYINPUT17), .Z(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n614_), .B2(new_n547_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n614_), .B2(new_n547_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n577_), .A2(new_n580_), .A3(new_n606_), .A4(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n516_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n424_), .B1(new_n423_), .B2(new_n341_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n340_), .A2(KEYINPUT100), .A3(new_n342_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n202_), .B1(new_n624_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n419_), .A2(new_n420_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n429_), .A2(new_n430_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n631_), .A2(new_n632_), .B1(new_n357_), .B2(new_n414_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n606_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n577_), .A2(new_n580_), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT37), .B1(new_n510_), .B2(new_n513_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT37), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n509_), .B(new_n638_), .C1(new_n504_), .C2(new_n512_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n636_), .A2(new_n641_), .A3(new_n621_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n635_), .A2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT101), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n202_), .A3(new_n628_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n646_));
  AOI21_X1  g445(.A(new_n629_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n646_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n644_), .A2(new_n202_), .A3(new_n648_), .A4(new_n628_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n647_), .B1(new_n651_), .B2(new_n652_), .ZN(G1324gat));
  XNOR2_X1  g452(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n633_), .A2(new_n514_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n623_), .A2(new_n421_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT104), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n432_), .A2(KEYINPUT104), .A3(new_n515_), .A4(new_n658_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G8gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n656_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n432_), .A2(new_n515_), .A3(new_n658_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n665_), .A2(KEYINPUT105), .A3(G8gat), .A4(new_n660_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n662_), .A2(KEYINPUT106), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT106), .B1(new_n662_), .B2(new_n666_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n662_), .A2(new_n666_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n669_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n630_), .A2(new_n581_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n644_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n655_), .B1(new_n670_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n671_), .A2(new_n672_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n662_), .A2(KEYINPUT106), .A3(new_n666_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(KEYINPUT39), .A3(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n680_), .A2(new_n673_), .A3(new_n675_), .A4(new_n654_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n677_), .A2(new_n681_), .ZN(G1325gat));
  AOI21_X1  g481(.A(new_n398_), .B1(new_n624_), .B2(new_n413_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT41), .ZN(new_n684_));
  INV_X1    g483(.A(new_n643_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n398_), .A3(new_n413_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1326gat));
  INV_X1    g486(.A(G22gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n624_), .B2(new_n396_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT42), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n685_), .A2(new_n688_), .A3(new_n396_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1327gat));
  NAND2_X1  g491(.A1(new_n514_), .A2(new_n621_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n636_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n635_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n628_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n432_), .A2(new_n641_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n622_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n636_), .A2(new_n634_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(KEYINPUT44), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n432_), .A2(KEYINPUT43), .A3(new_n641_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n699_), .A2(new_n700_), .A3(new_n703_), .A4(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n633_), .B2(new_n640_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n706_), .A2(new_n704_), .A3(new_n621_), .A4(new_n700_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n702_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n628_), .A2(G29gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n696_), .B1(new_n709_), .B2(new_n710_), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n705_), .A2(new_n708_), .A3(new_n630_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G36gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n421_), .A2(G36gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n635_), .A2(new_n694_), .A3(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT45), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT46), .B1(new_n717_), .B2(KEYINPUT109), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n719_), .B(new_n720_), .C1(new_n713_), .C2(new_n716_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1329gat));
  NAND3_X1  g521(.A1(new_n709_), .A2(G43gat), .A3(new_n413_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n695_), .A2(new_n413_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n406_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n723_), .A2(KEYINPUT47), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT47), .B1(new_n723_), .B2(new_n725_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n695_), .B2(new_n396_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n396_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n709_), .B2(new_n730_), .ZN(G1331gat));
  AOI21_X1  g530(.A(new_n621_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n432_), .A2(new_n634_), .A3(new_n732_), .A4(new_n636_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT110), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n628_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n519_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n736_), .A2(KEYINPUT111), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(KEYINPUT111), .ZN(new_n738_));
  INV_X1    g537(.A(new_n636_), .ZN(new_n739_));
  NOR4_X1   g538(.A1(new_n516_), .A2(new_n606_), .A3(new_n621_), .A4(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n627_), .A2(new_n519_), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n737_), .A2(new_n738_), .B1(new_n740_), .B2(new_n741_), .ZN(G1332gat));
  AOI21_X1  g541(.A(new_n517_), .B1(new_n740_), .B2(new_n630_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n630_), .A2(new_n517_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT113), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n734_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1333gat));
  NAND3_X1  g548(.A1(new_n734_), .A2(new_n524_), .A3(new_n413_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n740_), .A2(new_n413_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G71gat), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT49), .B(new_n524_), .C1(new_n740_), .C2(new_n413_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT114), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n740_), .A2(new_n396_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G78gat), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT115), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n758_), .B(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT50), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n734_), .A2(new_n526_), .A3(new_n396_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n764_), .A3(new_n765_), .ZN(G1335gat));
  NAND4_X1  g565(.A1(new_n699_), .A2(new_n634_), .A3(new_n636_), .A4(new_n704_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n767_), .A2(new_n627_), .A3(new_n452_), .ZN(new_n768_));
  NOR4_X1   g567(.A1(new_n633_), .A2(new_n606_), .A3(new_n739_), .A4(new_n693_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G85gat), .B1(new_n769_), .B2(new_n628_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1336gat));
  AOI21_X1  g570(.A(G92gat), .B1(new_n769_), .B2(new_n630_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT116), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n767_), .A2(new_n456_), .A3(new_n421_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1337gat));
  OAI21_X1  g574(.A(G99gat), .B1(new_n767_), .B2(new_n428_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n769_), .A2(new_n413_), .A3(new_n441_), .A4(new_n443_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n776_), .A2(new_n777_), .B1(KEYINPUT117), .B2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(KEYINPUT117), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(G1338gat));
  NAND3_X1  g580(.A1(new_n769_), .A2(new_n442_), .A3(new_n396_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT118), .ZN(new_n783_));
  INV_X1    g582(.A(new_n396_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G106gat), .B1(new_n767_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n786_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT53), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n785_), .A2(new_n786_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n788_), .A4(new_n783_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1339gat));
  INV_X1    g593(.A(new_n430_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n627_), .A2(new_n630_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  AND4_X1   g596(.A1(new_n560_), .A2(new_n551_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n551_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n562_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(KEYINPUT55), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n799_), .A2(new_n802_), .A3(new_n562_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n797_), .B(new_n570_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n592_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n594_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n589_), .A2(new_n591_), .A3(new_n805_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  MUX2_X1   g607(.A(new_n808_), .B(new_n595_), .S(new_n603_), .Z(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(new_n573_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n804_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n570_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT58), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT120), .B1(new_n814_), .B2(new_n640_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n811_), .A2(KEYINPUT58), .A3(new_n813_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n802_), .B1(new_n799_), .B2(new_n562_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(new_n798_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n797_), .B1(new_n819_), .B2(new_n570_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n804_), .A2(new_n810_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n817_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n641_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n815_), .A2(new_n816_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NOR2_X1   g625(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n812_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n570_), .B(new_n827_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n606_), .A2(new_n573_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n809_), .B1(new_n579_), .B2(new_n574_), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n826_), .B(new_n514_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n827_), .B1(new_n819_), .B2(new_n570_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n830_), .A2(new_n831_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT57), .B1(new_n837_), .B2(new_n515_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n834_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n622_), .B1(new_n825_), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n739_), .A2(new_n634_), .A3(new_n732_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n795_), .B(new_n796_), .C1(new_n840_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(G113gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n606_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n824_), .A2(new_n816_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n823_), .B1(new_n822_), .B2(new_n641_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n838_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n837_), .A2(KEYINPUT57), .A3(new_n515_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n621_), .B1(new_n850_), .B2(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n841_), .B(KEYINPUT54), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n856_), .A2(KEYINPUT59), .A3(new_n795_), .A4(new_n796_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n844_), .A2(new_n858_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n857_), .A2(new_n859_), .A3(KEYINPUT121), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT121), .B1(new_n857_), .B2(new_n859_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n634_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n847_), .B1(new_n862_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g662(.A(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n739_), .B2(KEYINPUT60), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n845_), .B(new_n865_), .C1(KEYINPUT60), .C2(new_n864_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n739_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n864_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n845_), .B2(new_n622_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n860_), .A2(new_n861_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n621_), .A2(KEYINPUT122), .ZN(new_n871_));
  MUX2_X1   g670(.A(KEYINPUT122), .B(new_n871_), .S(G127gat), .Z(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n870_), .B2(new_n872_), .ZN(G1342gat));
  AOI21_X1  g672(.A(G134gat), .B1(new_n845_), .B2(new_n514_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n641_), .A2(G134gat), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT123), .Z(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n870_), .B2(new_n876_), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n840_), .A2(new_n843_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n627_), .A2(new_n429_), .A3(new_n630_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT124), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n606_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n636_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n622_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1346gat));
  INV_X1    g687(.A(G162gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n881_), .A2(new_n889_), .A3(new_n514_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n881_), .A2(new_n641_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n892_), .B2(new_n889_), .ZN(G1347gat));
  XNOR2_X1  g692(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n627_), .A2(new_n630_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n856_), .A2(new_n795_), .A3(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n634_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT22), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n894_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(G169gat), .ZN(new_n901_));
  INV_X1    g700(.A(G169gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n898_), .B2(new_n894_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n900_), .B2(new_n903_), .ZN(G1348gat));
  NOR2_X1   g703(.A1(new_n897_), .A2(new_n739_), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(G176gat), .Z(G1349gat));
  NOR2_X1   g705(.A1(new_n897_), .A2(new_n621_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(G183gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n258_), .B2(new_n907_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n897_), .B2(new_n640_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n515_), .A2(new_n259_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n897_), .B2(new_n911_), .ZN(G1351gat));
  NOR3_X1   g711(.A1(new_n878_), .A2(new_n429_), .A3(new_n895_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n606_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT126), .B(G197gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1352gat));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n636_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g717(.A1(new_n913_), .A2(new_n622_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  NAND2_X1  g722(.A1(new_n913_), .A2(new_n641_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G218gat), .ZN(new_n925_));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n913_), .A2(new_n926_), .A3(new_n514_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n925_), .A2(KEYINPUT127), .A3(new_n927_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1355gat));
endmodule


