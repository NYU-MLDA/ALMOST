//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT68), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n210_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT66), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  INV_X1    g023(.A(G92gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n220_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n219_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n208_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT65), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n217_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n223_), .A2(new_n228_), .A3(new_n237_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n236_), .A2(KEYINPUT67), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT67), .B1(new_n236_), .B2(new_n238_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n232_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  OAI22_X1  g040(.A1(new_n221_), .A2(new_n222_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n243_));
  XOR2_X1   g042(.A(KEYINPUT10), .B(G99gat), .Z(new_n244_));
  AOI22_X1  g043(.A1(new_n242_), .A2(new_n243_), .B1(new_n244_), .B2(new_n213_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n242_), .A2(new_n243_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT65), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT65), .B1(new_n205_), .B2(new_n207_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G29gat), .B(G36gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT72), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n252_), .A2(new_n253_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G43gat), .B(G50gat), .Z(new_n256_));
  OR3_X1    g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n203_), .B1(new_n251_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n250_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n247_), .A2(new_n248_), .A3(new_n216_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n223_), .A2(new_n228_), .A3(new_n237_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n236_), .A2(new_n238_), .A3(KEYINPUT67), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n261_), .B1(new_n267_), .B2(new_n232_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n259_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(KEYINPUT74), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n260_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n237_), .B1(new_n219_), .B2(new_n230_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n274_), .B2(new_n261_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n241_), .A2(KEYINPUT71), .A3(new_n250_), .ZN(new_n276_));
  XOR2_X1   g075(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n259_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n259_), .A2(new_n278_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n275_), .B(new_n276_), .C1(new_n279_), .C2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G232gat), .A2(G233gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT34), .Z(new_n284_));
  INV_X1    g083(.A(KEYINPUT35), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n286_), .B(KEYINPUT75), .Z(new_n287_));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n271_), .A2(new_n282_), .A3(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n284_), .A2(new_n285_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n289_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n260_), .B2(new_n270_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n291_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n282_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G190gat), .B(G218gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT76), .ZN(new_n298_));
  XOR2_X1   g097(.A(G134gat), .B(G162gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(KEYINPUT36), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n292_), .A2(new_n296_), .A3(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n300_), .B(KEYINPUT36), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n303_), .A2(new_n306_), .A3(KEYINPUT37), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT37), .ZN(new_n308_));
  INV_X1    g107(.A(new_n296_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n295_), .B1(new_n294_), .B2(new_n282_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n304_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n292_), .A2(new_n296_), .A3(new_n302_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n308_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n307_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G127gat), .B(G155gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G183gat), .B(G211gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT17), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G15gat), .B(G22gat), .ZN(new_n321_));
  INV_X1    g120(.A(G1gat), .ZN(new_n322_));
  INV_X1    g121(.A(G8gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT14), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G1gat), .B(G8gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  NAND2_X1  g126(.A1(G231gat), .A2(G233gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n328_), .B(KEYINPUT78), .Z(new_n329_));
  XOR2_X1   g128(.A(new_n327_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G57gat), .B(G64gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT11), .ZN(new_n333_));
  XOR2_X1   g132(.A(G71gat), .B(G78gat), .Z(new_n334_));
  OR2_X1    g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n334_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n332_), .A2(KEYINPUT11), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT69), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n320_), .B1(new_n331_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n331_), .B2(new_n339_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n319_), .A2(KEYINPUT17), .ZN(new_n342_));
  INV_X1    g141(.A(new_n338_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n330_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n343_), .B2(new_n330_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n314_), .A2(KEYINPUT80), .A3(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT80), .B1(new_n314_), .B2(new_n347_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OR4_X1    g149(.A1(KEYINPUT90), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n351_));
  OR2_X1    g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT3), .B1(new_n352_), .B2(KEYINPUT90), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G141gat), .A2(G148gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT87), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT2), .ZN(new_n357_));
  NAND3_X1  g156(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n351_), .A2(new_n353_), .A3(new_n359_), .A4(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G155gat), .ZN(new_n362_));
  INV_X1    g161(.A(G162gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT88), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT88), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(G155gat), .B2(G162gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n367_), .B1(G155gat), .B2(G162gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n361_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT97), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT1), .B1(new_n362_), .B2(new_n363_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT1), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(G155gat), .A3(G162gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n371_), .A2(new_n364_), .A3(new_n366_), .A4(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n356_), .A2(new_n352_), .A3(new_n358_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(KEYINPUT89), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT89), .B1(new_n374_), .B2(new_n375_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n369_), .B(new_n370_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G127gat), .B(G134gat), .Z(new_n380_));
  XOR2_X1   g179(.A(G113gat), .B(G120gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n374_), .A2(new_n375_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT89), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n376_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n382_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n370_), .A4(new_n369_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT4), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n369_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n382_), .A2(KEYINPUT4), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n391_), .A2(new_n398_), .A3(KEYINPUT98), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT98), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n383_), .B2(new_n389_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n402_), .B2(new_n397_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n390_), .A2(new_n395_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(G85gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT0), .B(G57gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n399_), .A2(new_n403_), .A3(new_n404_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n408_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n390_), .B2(new_n396_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n394_), .A2(new_n395_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n402_), .B2(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT96), .ZN(new_n417_));
  INV_X1    g216(.A(G197gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT91), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G197gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n421_), .A3(G204gat), .ZN(new_n422_));
  INV_X1    g221(.A(G204gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT93), .B1(new_n423_), .B2(G197gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT91), .B(G197gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT94), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n425_), .A2(new_n427_), .A3(KEYINPUT94), .ZN(new_n431_));
  XOR2_X1   g230(.A(G211gat), .B(G218gat), .Z(new_n432_));
  AND2_X1   g231(.A1(new_n432_), .A2(KEYINPUT21), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT21), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n418_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT92), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n423_), .B2(G197gat), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n437_), .B(new_n439_), .C1(new_n426_), .C2(G204gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n432_), .B1(new_n440_), .B2(KEYINPUT21), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n434_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT23), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G169gat), .ZN(new_n449_));
  INV_X1    g248(.A(G176gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(KEYINPUT24), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G169gat), .A2(G176gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(KEYINPUT24), .A3(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n448_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT25), .B(G183gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT26), .B(G190gat), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n446_), .B(new_n447_), .C1(G183gat), .C2(G190gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT22), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n443_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G190gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT83), .B1(new_n467_), .B2(KEYINPUT26), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n456_), .B(new_n468_), .C1(new_n457_), .C2(KEYINPUT83), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n464_), .B1(new_n470_), .B2(new_n455_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT84), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n469_), .A2(new_n448_), .A3(new_n454_), .A4(new_n452_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n464_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n472_), .A2(new_n442_), .A3(new_n434_), .A4(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n466_), .A2(new_n476_), .A3(KEYINPUT20), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G226gat), .A2(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT19), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G8gat), .B(G36gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(G64gat), .B(G92gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n475_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n474_), .B1(new_n473_), .B2(new_n464_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n443_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n479_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n434_), .A2(new_n442_), .A3(new_n464_), .A4(new_n459_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n489_), .A2(KEYINPUT20), .A3(new_n490_), .A4(new_n491_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n480_), .A2(new_n486_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n486_), .B1(new_n480_), .B2(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n417_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n399_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n409_), .B1(new_n496_), .B2(new_n408_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n480_), .A2(new_n492_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n485_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n480_), .A2(new_n486_), .A3(new_n492_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(KEYINPUT96), .A3(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n416_), .A2(new_n495_), .A3(new_n497_), .A4(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n477_), .A2(new_n479_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n491_), .A2(KEYINPUT20), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n472_), .A2(new_n475_), .B1(new_n434_), .B2(new_n442_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n479_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT99), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT99), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n508_), .B(new_n479_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n503_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n486_), .A2(KEYINPUT32), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n498_), .A2(new_n511_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n496_), .A2(new_n408_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n402_), .A2(new_n397_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n515_), .A2(KEYINPUT98), .B1(new_n390_), .B2(new_n395_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n412_), .B1(new_n516_), .B2(new_n403_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n512_), .B(new_n513_), .C1(new_n514_), .C2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n502_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G227gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(G15gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G71gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n521_), .B(G15gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(G71gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n212_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(G71gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(new_n524_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(G99gat), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT85), .B(G43gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT30), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n528_), .A2(new_n531_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n472_), .A2(new_n536_), .A3(new_n475_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n535_), .B1(new_n533_), .B2(new_n537_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n520_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n537_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n535_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(KEYINPUT86), .A3(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n382_), .B(KEYINPUT31), .Z(new_n546_));
  NAND3_X1  g345(.A1(new_n540_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n520_), .B(new_n548_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G228gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(G78gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(new_n213_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G22gat), .B(G50gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT28), .B1(new_n392_), .B2(KEYINPUT29), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n386_), .A2(new_n376_), .B1(new_n361_), .B2(new_n368_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT28), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n392_), .A2(KEYINPUT29), .B1(new_n442_), .B2(new_n434_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n443_), .B1(new_n562_), .B2(new_n560_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n559_), .B2(new_n563_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n558_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n565_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n557_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n551_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n519_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n550_), .A2(new_n573_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n569_), .A2(new_n572_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n510_), .A2(new_n485_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n493_), .A2(KEYINPUT100), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n500_), .A2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n583_), .A2(new_n584_), .A3(KEYINPUT27), .A4(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n514_), .A2(new_n517_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n579_), .A2(new_n582_), .A3(new_n587_), .A4(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n575_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT70), .B1(new_n251_), .B2(new_n339_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT70), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT69), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n338_), .B(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n268_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n268_), .A2(new_n595_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n591_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n343_), .A2(KEYINPUT12), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n275_), .A2(new_n276_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n268_), .B2(new_n595_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n591_), .B1(new_n268_), .B2(new_n595_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n602_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT5), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n599_), .A2(new_n606_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n599_), .B2(new_n606_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT13), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT13), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G113gat), .B(G141gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT81), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n269_), .A2(new_n277_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n327_), .B1(new_n626_), .B2(new_n280_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n327_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n259_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n627_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n631_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n259_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n628_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n625_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n630_), .B1(new_n281_), .B2(new_n279_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n628_), .A3(new_n633_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n635_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n624_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n636_), .A2(KEYINPUT82), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT82), .B1(new_n636_), .B2(new_n640_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n590_), .A2(new_n620_), .A3(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n350_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n588_), .B(KEYINPUT102), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(G1gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(KEYINPUT103), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650_));
  INV_X1    g449(.A(new_n644_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n349_), .A3(new_n348_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n647_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n648_), .A2(new_n649_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n649_), .B1(new_n648_), .B2(new_n654_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n202_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n648_), .A2(new_n654_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT104), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(KEYINPUT38), .A3(new_n655_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n588_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n587_), .A2(new_n582_), .ZN(new_n664_));
  AOI22_X1  g463(.A1(new_n663_), .A2(new_n664_), .B1(new_n519_), .B2(new_n574_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n311_), .A2(new_n312_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n643_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n619_), .A2(new_n347_), .A3(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G1gat), .B1(new_n672_), .B2(new_n588_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n658_), .A2(new_n661_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT105), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n658_), .A2(new_n661_), .A3(new_n676_), .A4(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1324gat));
  INV_X1    g477(.A(new_n664_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n671_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G8gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT39), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n645_), .A2(new_n323_), .A3(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1325gat));
  NAND3_X1  g485(.A1(new_n645_), .A2(new_n522_), .A3(new_n551_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n671_), .A2(new_n551_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n688_), .B2(G15gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT107), .Z(G1326gat));
  INV_X1    g491(.A(G22gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n671_), .B2(new_n573_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT42), .Z(new_n695_));
  NAND3_X1  g494(.A1(new_n645_), .A2(new_n693_), .A3(new_n573_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1327gat));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  INV_X1    g497(.A(new_n314_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n665_), .A2(new_n699_), .A3(KEYINPUT43), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(new_n307_), .B2(new_n313_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT37), .B1(new_n303_), .B2(new_n306_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n311_), .A2(new_n308_), .A3(new_n312_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(KEYINPUT108), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n706_), .B2(new_n665_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT109), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n590_), .A2(new_n702_), .A3(new_n705_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(KEYINPUT43), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n700_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n619_), .A2(new_n669_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n347_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n698_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n700_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n709_), .A2(new_n710_), .A3(KEYINPUT43), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n710_), .B1(new_n709_), .B2(KEYINPUT43), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n719_), .A2(KEYINPUT44), .A3(new_n347_), .A4(new_n713_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n646_), .ZN(new_n721_));
  AND4_X1   g520(.A1(G29gat), .A2(new_n715_), .A3(new_n720_), .A4(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n666_), .A2(new_n346_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT110), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n724_), .A2(new_n620_), .A3(new_n590_), .A4(new_n643_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT111), .ZN(new_n726_));
  AOI21_X1  g525(.A(G29gat), .B1(new_n726_), .B2(new_n662_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n722_), .A2(new_n727_), .ZN(G1328gat));
  INV_X1    g527(.A(new_n726_), .ZN(new_n729_));
  INV_X1    g528(.A(G36gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n679_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT45), .B1(new_n729_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n726_), .A2(new_n733_), .A3(new_n730_), .A4(new_n679_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n715_), .A2(new_n720_), .A3(new_n679_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G36gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n737_), .A3(KEYINPUT46), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1329gat));
  NAND4_X1  g541(.A1(new_n715_), .A2(new_n720_), .A3(G43gat), .A4(new_n551_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n729_), .A2(new_n550_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(G43gat), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g545(.A1(new_n715_), .A2(new_n720_), .A3(new_n573_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G50gat), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n577_), .A2(G50gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n726_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n748_), .A2(KEYINPUT113), .A3(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1331gat));
  NAND4_X1  g555(.A1(new_n668_), .A2(new_n346_), .A3(new_n619_), .A4(new_n669_), .ZN(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n588_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n665_), .A2(new_n643_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n619_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(new_n350_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n646_), .B1(new_n763_), .B2(KEYINPUT114), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(KEYINPUT114), .B2(new_n763_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n759_), .B1(new_n765_), .B2(new_n758_), .ZN(G1332gat));
  OAI21_X1  g565(.A(G64gat), .B1(new_n757_), .B2(new_n664_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT48), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n664_), .A2(G64gat), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT115), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(new_n763_), .B2(new_n770_), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n757_), .B2(new_n550_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n762_), .A2(new_n524_), .A3(new_n551_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1334gat));
  OAI21_X1  g575(.A(G78gat), .B1(new_n757_), .B2(new_n577_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT50), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n573_), .A2(new_n553_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT117), .Z(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n763_), .B2(new_n780_), .ZN(G1335gat));
  AND3_X1   g580(.A1(new_n760_), .A2(new_n619_), .A3(new_n724_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n224_), .A3(new_n721_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n619_), .A2(new_n347_), .A3(new_n669_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n712_), .A2(new_n588_), .A3(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n785_), .B2(new_n224_), .ZN(G1336gat));
  NOR2_X1   g585(.A1(new_n712_), .A2(new_n784_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n225_), .B1(new_n787_), .B2(new_n679_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n664_), .A2(G92gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n782_), .B2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT118), .ZN(G1337gat));
  AOI21_X1  g590(.A(new_n212_), .B1(new_n787_), .B2(new_n551_), .ZN(new_n792_));
  AND2_X1   g591(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n782_), .A2(new_n244_), .A3(new_n551_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(G1338gat));
  INV_X1    g596(.A(new_n784_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n719_), .A2(new_n573_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(new_n800_), .A3(G106gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n799_), .B2(G106gat), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n712_), .A2(new_n577_), .A3(new_n784_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT120), .B(new_n803_), .C1(new_n805_), .C2(new_n213_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n577_), .A2(G106gat), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n782_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT53), .B1(new_n804_), .B2(new_n809_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n802_), .A2(new_n803_), .B1(new_n782_), .B2(new_n807_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT120), .B1(new_n805_), .B2(new_n213_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT52), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n811_), .B(new_n812_), .C1(new_n814_), .C2(new_n801_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n810_), .A2(new_n815_), .ZN(G1339gat));
  NOR4_X1   g615(.A1(new_n314_), .A2(new_n619_), .A3(new_n347_), .A4(new_n643_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT54), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n627_), .A2(new_n631_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n819_), .A2(KEYINPUT122), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(KEYINPUT122), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n629_), .A3(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n633_), .A2(new_n634_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n822_), .B(new_n625_), .C1(new_n629_), .C2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n640_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n613_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n606_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n606_), .A2(KEYINPUT121), .A3(new_n827_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n602_), .A2(new_n604_), .A3(new_n605_), .A4(KEYINPUT55), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n602_), .A2(new_n604_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n591_), .B1(new_n833_), .B2(new_n597_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .A4(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n835_), .B2(new_n610_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(KEYINPUT123), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n839_));
  AOI211_X1 g638(.A(new_n839_), .B(KEYINPUT56), .C1(new_n835_), .C2(new_n610_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT58), .B(new_n826_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n826_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n699_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n845_), .B2(KEYINPUT124), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n835_), .A2(new_n610_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n839_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n837_), .A2(KEYINPUT123), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n836_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT58), .B1(new_n853_), .B2(new_n826_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n847_), .B1(new_n854_), .B2(new_n699_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n846_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n643_), .A2(new_n612_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n850_), .B2(new_n836_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n825_), .A2(new_n615_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n666_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT57), .B(new_n666_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n856_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n818_), .B1(new_n866_), .B2(new_n347_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n646_), .A2(new_n679_), .A3(new_n578_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT125), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G113gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n818_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n864_), .B1(new_n846_), .B2(new_n855_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n346_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n868_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n870_), .A2(new_n871_), .A3(new_n643_), .A4(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n874_), .A2(KEYINPUT59), .A3(new_n868_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n669_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n877_), .B1(new_n881_), .B2(new_n871_), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n883_), .A2(KEYINPUT60), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n620_), .B2(KEYINPUT60), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n870_), .A2(new_n876_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n620_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n883_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n870_), .A2(new_n889_), .A3(new_n346_), .A4(new_n876_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n347_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1342gat));
  INV_X1    g691(.A(G134gat), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n870_), .A2(new_n893_), .A3(new_n667_), .A4(new_n876_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n699_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n893_), .ZN(G1343gat));
  NOR3_X1   g695(.A1(new_n646_), .A2(new_n679_), .A3(new_n576_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n874_), .A2(new_n643_), .A3(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT126), .B(G141gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1344gat));
  INV_X1    g699(.A(new_n897_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n867_), .A2(new_n620_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(G148gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1345gat));
  NOR3_X1   g703(.A1(new_n867_), .A2(new_n347_), .A3(new_n901_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT61), .B(G155gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1346gat));
  NOR2_X1   g706(.A1(new_n867_), .A2(new_n901_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G162gat), .B1(new_n908_), .B2(new_n667_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n706_), .A2(new_n363_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n908_), .B2(new_n910_), .ZN(G1347gat));
  NOR3_X1   g710(.A1(new_n721_), .A2(new_n664_), .A3(new_n550_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n912_), .A2(new_n643_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n874_), .A2(new_n462_), .A3(new_n577_), .A4(new_n913_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n914_), .A2(KEYINPUT62), .A3(new_n449_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(KEYINPUT62), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n874_), .A2(new_n917_), .A3(new_n577_), .A4(new_n913_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n918_), .A2(G169gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n915_), .B1(new_n916_), .B2(new_n919_), .ZN(G1348gat));
  NAND4_X1  g719(.A1(new_n874_), .A2(new_n619_), .A3(new_n577_), .A4(new_n912_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g721(.A1(new_n874_), .A2(new_n346_), .A3(new_n577_), .A4(new_n912_), .ZN(new_n923_));
  MUX2_X1   g722(.A(new_n456_), .B(G183gat), .S(new_n923_), .Z(G1350gat));
  NOR2_X1   g723(.A1(new_n867_), .A2(new_n573_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n925_), .A2(new_n667_), .A3(new_n457_), .A4(new_n912_), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n925_), .A2(new_n314_), .A3(new_n912_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n467_), .ZN(G1351gat));
  NOR3_X1   g727(.A1(new_n664_), .A2(new_n662_), .A3(new_n576_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n874_), .A2(new_n643_), .A3(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n620_), .B1(new_n932_), .B2(G204gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n874_), .A2(new_n929_), .A3(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n423_), .A2(KEYINPUT127), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n874_), .A2(new_n346_), .A3(new_n929_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  AND2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n937_), .A2(new_n938_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n940_), .B1(new_n937_), .B2(new_n938_), .ZN(G1354gat));
  INV_X1    g740(.A(G218gat), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n874_), .A2(new_n942_), .A3(new_n667_), .A4(new_n929_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n929_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n867_), .A2(new_n699_), .A3(new_n944_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n945_), .B2(new_n942_), .ZN(G1355gat));
endmodule


