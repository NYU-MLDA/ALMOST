//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_;
  INV_X1    g000(.A(G92gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT65), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G92gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n205_), .A3(G85gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(new_n202_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n211_), .B1(new_n213_), .B2(KEYINPUT9), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n206_), .A2(KEYINPUT66), .A3(new_n207_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n210_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT10), .B(G99gat), .Z(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n216_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n213_), .A2(new_n211_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n219_), .B(new_n220_), .C1(new_n227_), .C2(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n229_), .B(new_n223_), .C1(new_n230_), .C2(KEYINPUT67), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n227_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n226_), .B1(new_n228_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT8), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n236_), .B(new_n226_), .C1(new_n228_), .C2(new_n233_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n225_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G29gat), .ZN(new_n240_));
  INV_X1    g039(.A(G36gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G43gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G29gat), .A2(G36gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G50gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G29gat), .B(G36gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G43gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(G50gat), .B1(new_n251_), .B2(new_n245_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT74), .B1(new_n239_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT74), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n225_), .A2(new_n238_), .A3(new_n256_), .A4(new_n253_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G232gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT71), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT34), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT73), .B1(new_n249_), .B2(new_n252_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n247_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n251_), .A2(G50gat), .A3(new_n245_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n266_), .A2(KEYINPUT15), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT15), .B1(new_n266_), .B2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n239_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n261_), .A2(new_n263_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n258_), .A2(new_n265_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n276_), .A2(KEYINPUT75), .A3(new_n264_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT75), .B1(new_n276_), .B2(new_n264_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n275_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G190gat), .B(G218gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G134gat), .ZN(new_n281_));
  INV_X1    g080(.A(G162gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(KEYINPUT36), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(KEYINPUT36), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n279_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT76), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n285_), .B(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n275_), .B(new_n289_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(KEYINPUT77), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT37), .ZN(new_n292_));
  INV_X1    g091(.A(new_n290_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n287_), .A2(new_n290_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT37), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n291_), .A2(new_n295_), .A3(KEYINPUT78), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G15gat), .B(G22gat), .ZN(new_n304_));
  INV_X1    g103(.A(G1gat), .ZN(new_n305_));
  INV_X1    g104(.A(G8gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT14), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G8gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G231gat), .A2(G233gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  XNOR2_X1  g111(.A(G57gat), .B(G64gat), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n313_), .A2(KEYINPUT11), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(KEYINPUT11), .ZN(new_n315_));
  XOR2_X1   g114(.A(G71gat), .B(G78gat), .Z(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n315_), .A2(new_n316_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n317_), .A2(KEYINPUT68), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT68), .B1(new_n317_), .B2(new_n318_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n312_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT16), .B(G183gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G211gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(G127gat), .B(G155gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT17), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n326_), .A2(new_n327_), .ZN(new_n329_));
  OR3_X1    g128(.A1(new_n322_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n317_), .A2(new_n318_), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n312_), .B(new_n331_), .Z(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n303_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT79), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G127gat), .A2(G134gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G127gat), .A2(G134gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(G113gat), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G127gat), .ZN(new_n342_));
  INV_X1    g141(.A(G134gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G113gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n338_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n341_), .A2(G120gat), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(G120gat), .B1(new_n341_), .B2(new_n346_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT83), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(KEYINPUT1), .ZN(new_n353_));
  OR2_X1    g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(KEYINPUT1), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n356_), .A2(KEYINPUT83), .A3(G155gat), .A4(G162gat), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .A4(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G141gat), .A2(G148gat), .ZN(new_n359_));
  INV_X1    g158(.A(G141gat), .ZN(new_n360_));
  INV_X1    g159(.A(G148gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n364_));
  NOR2_X1   g163(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n362_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n359_), .A2(KEYINPUT2), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT2), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(G141gat), .A3(G148gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n366_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT85), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n366_), .A2(new_n370_), .A3(new_n375_), .A4(new_n372_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n354_), .A2(new_n352_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n350_), .B(new_n363_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n349_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(KEYINPUT82), .A3(new_n347_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n378_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n363_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n381_), .B(new_n383_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n379_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n379_), .A2(new_n386_), .A3(KEYINPUT4), .ZN(new_n389_));
  INV_X1    g188(.A(new_n387_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n386_), .B2(KEYINPUT4), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n388_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n388_), .B(new_n397_), .C1(new_n389_), .C2(new_n391_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(KEYINPUT94), .A3(new_n398_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G22gat), .B(G50gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT28), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT29), .B1(new_n384_), .B2(new_n385_), .ZN(new_n408_));
  AND2_X1   g207(.A1(G211gat), .A2(G218gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G211gat), .A2(G218gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(G204gat), .ZN(new_n412_));
  AND2_X1   g211(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT21), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(G197gat), .B2(G204gat), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n411_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(G204gat), .B1(new_n413_), .B2(new_n414_), .ZN(new_n419_));
  INV_X1    g218(.A(G197gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(G204gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n416_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n422_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(KEYINPUT21), .A3(new_n411_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n408_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G228gat), .ZN(new_n429_));
  INV_X1    g228(.A(G233gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n408_), .B(new_n427_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT86), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT29), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n436_), .B(new_n363_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n432_), .A2(new_n441_), .A3(new_n433_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n435_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n440_), .B1(new_n435_), .B2(new_n442_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n407_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n406_), .A3(new_n443_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G169gat), .A2(G176gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT24), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT88), .ZN(new_n452_));
  INV_X1    g251(.A(G169gat), .ZN(new_n453_));
  INV_X1    g252(.A(G176gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n450_), .A2(new_n456_), .A3(KEYINPUT24), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n452_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT24), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G183gat), .A2(G190gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT23), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n460_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT25), .B(G183gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n458_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(G183gat), .A2(G190gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n463_), .A2(new_n472_), .A3(new_n464_), .ZN(new_n473_));
  AND2_X1   g272(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n454_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n473_), .A2(new_n476_), .A3(new_n450_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n424_), .A2(new_n471_), .A3(new_n426_), .A4(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n477_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT25), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G183gat), .ZN(new_n481_));
  INV_X1    g280(.A(G183gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT25), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT81), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT81), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n466_), .A2(new_n467_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n451_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n485_), .A2(new_n487_), .B1(new_n455_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n479_), .B1(new_n489_), .B2(new_n465_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n411_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n492_), .A2(KEYINPUT21), .B1(new_n418_), .B2(new_n423_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n478_), .B(KEYINPUT20), .C1(new_n490_), .C2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G226gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT19), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n471_), .A2(new_n477_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n427_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n496_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n488_), .A2(new_n455_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n481_), .A2(new_n486_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n468_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n486_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n465_), .B(new_n501_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n505_), .A2(new_n424_), .A3(new_n426_), .A4(new_n477_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n499_), .A2(KEYINPUT20), .A3(new_n500_), .A4(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n497_), .A2(KEYINPUT92), .A3(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n507_), .A2(KEYINPUT92), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G8gat), .B(G36gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G64gat), .B(G92gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT96), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n515_), .A2(KEYINPUT96), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n508_), .A2(new_n509_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n499_), .A2(KEYINPUT20), .A3(new_n496_), .A4(new_n506_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n505_), .A2(new_n477_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n522_), .B2(new_n427_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n496_), .B1(new_n523_), .B2(new_n478_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n514_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n518_), .A2(KEYINPUT27), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n494_), .A2(new_n500_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(new_n515_), .A3(new_n519_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT98), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT98), .ZN(new_n533_));
  AOI211_X1 g332(.A(new_n533_), .B(new_n530_), .C1(new_n525_), .C2(new_n528_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n526_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT99), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n526_), .B(KEYINPUT99), .C1(new_n532_), .C2(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n383_), .A2(new_n381_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n540_), .B1(new_n383_), .B2(new_n381_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n542_), .A2(new_n522_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n522_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G15gat), .B(G43gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT31), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n545_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G71gat), .B(G99gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G227gat), .A2(G233gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  AND2_X1   g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n552_), .A2(new_n555_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AND4_X1   g357(.A1(new_n404_), .A2(new_n449_), .A3(new_n539_), .A4(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n520_), .A2(new_n524_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n514_), .A2(KEYINPUT32), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n507_), .A2(KEYINPUT92), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n507_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT93), .B1(new_n568_), .B2(new_n562_), .ZN(new_n569_));
  AND4_X1   g368(.A1(KEYINPUT93), .A2(new_n508_), .A3(new_n509_), .A4(new_n562_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n564_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n560_), .B1(new_n404_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n401_), .A2(KEYINPUT91), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT33), .ZN(new_n574_));
  INV_X1    g373(.A(new_n529_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n379_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n387_), .B1(new_n386_), .B2(KEYINPUT4), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n398_), .B(new_n576_), .C1(new_n389_), .C2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n401_), .A2(KEYINPUT91), .A3(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n574_), .A2(new_n575_), .A3(new_n578_), .A4(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n508_), .A2(new_n509_), .A3(new_n562_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n568_), .A2(KEYINPUT93), .A3(new_n562_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n563_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n586_), .A2(KEYINPUT95), .A3(new_n403_), .A4(new_n402_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n572_), .A2(new_n581_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n449_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n446_), .A2(new_n448_), .B1(new_n403_), .B2(new_n402_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n535_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n558_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n559_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n310_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n254_), .A2(new_n310_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n253_), .B(new_n310_), .Z(new_n600_));
  INV_X1    g399(.A(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G113gat), .B(G141gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n453_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(new_n420_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n599_), .A2(new_n602_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT80), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n599_), .A2(new_n602_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n605_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT13), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(new_n412_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT5), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n454_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n225_), .A2(new_n238_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n618_), .B1(new_n619_), .B2(new_n321_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT64), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n321_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT12), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n225_), .B2(new_n238_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n331_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n620_), .A2(new_n623_), .A3(new_n624_), .A4(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT70), .ZN(new_n629_));
  AOI22_X1  g428(.A1(new_n619_), .A2(new_n321_), .B1(new_n626_), .B2(new_n331_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT70), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n623_), .A4(new_n620_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n619_), .B(new_n321_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n622_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n617_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n635_), .A3(new_n617_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n613_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n640_), .A2(KEYINPUT13), .A3(new_n636_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n612_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n595_), .A2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n337_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n404_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n305_), .A3(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT38), .ZN(new_n647_));
  INV_X1    g446(.A(new_n299_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n595_), .A2(new_n648_), .A3(new_n334_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n642_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n642_), .A2(new_n650_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n654_), .B2(new_n404_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n647_), .A2(new_n655_), .ZN(G1324gat));
  INV_X1    g455(.A(new_n539_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n644_), .A2(new_n306_), .A3(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT101), .ZN(new_n659_));
  OAI21_X1  g458(.A(G8gat), .B1(new_n654_), .B2(new_n539_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT39), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n654_), .B2(new_n594_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  INV_X1    g464(.A(G15gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n644_), .A2(new_n666_), .A3(new_n558_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n654_), .B2(new_n449_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT42), .ZN(new_n670_));
  INV_X1    g469(.A(G22gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n449_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n644_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT102), .Z(G1327gat));
  INV_X1    g474(.A(new_n653_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n335_), .B1(new_n676_), .B2(new_n651_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n449_), .A2(new_n539_), .A3(new_n404_), .A4(new_n558_), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n588_), .A2(new_n449_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(new_n558_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n291_), .A2(new_n295_), .A3(KEYINPUT78), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT78), .B1(new_n291_), .B2(new_n295_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n300_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n680_), .A2(new_n681_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n681_), .B1(new_n680_), .B2(new_n684_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n677_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n595_), .B2(new_n303_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n680_), .A2(new_n684_), .A3(new_n681_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n692_), .A2(KEYINPUT103), .A3(KEYINPUT44), .A4(new_n677_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n677_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n689_), .A2(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(new_n645_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n299_), .A2(new_n335_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n643_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n645_), .A2(new_n240_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT104), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n697_), .A2(new_n240_), .B1(new_n700_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n689_), .A2(new_n693_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n539_), .B1(new_n695_), .B2(new_n694_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n241_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n643_), .A2(new_n657_), .A3(new_n698_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n709_));
  OR3_X1    g508(.A1(new_n708_), .A2(G36gat), .A3(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G36gat), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n704_), .B1(new_n707_), .B2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n710_), .A2(new_n711_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n334_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n657_), .B1(new_n716_), .B2(KEYINPUT44), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT106), .B(new_n714_), .C1(new_n718_), .C2(new_n241_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n713_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT107), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n713_), .A2(new_n719_), .A3(new_n723_), .A4(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n707_), .A2(new_n720_), .A3(new_n712_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT108), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1329gat));
  OAI21_X1  g527(.A(new_n243_), .B1(new_n700_), .B2(new_n594_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n594_), .A2(new_n243_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n696_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n696_), .B2(new_n731_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g534(.A(G50gat), .B1(new_n699_), .B2(new_n672_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n449_), .A2(new_n247_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n696_), .B2(new_n737_), .ZN(G1331gat));
  OR2_X1    g537(.A1(new_n639_), .A2(new_n641_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(new_n612_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n649_), .A2(G57gat), .A3(new_n645_), .A4(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n680_), .A2(new_n740_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n337_), .A2(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n404_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n741_), .B1(new_n744_), .B2(G57gat), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT110), .Z(G1332gat));
  NAND2_X1  g545(.A1(new_n649_), .A2(new_n740_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G64gat), .B1(new_n747_), .B2(new_n539_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT48), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n539_), .A2(G64gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n743_), .B2(new_n750_), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n747_), .B2(new_n594_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT49), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n743_), .A2(G71gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n594_), .ZN(G1334gat));
  OAI21_X1  g554(.A(G78gat), .B1(new_n747_), .B2(new_n449_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n449_), .A2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n743_), .B2(new_n758_), .ZN(G1335gat));
  NAND2_X1  g558(.A1(new_n742_), .A2(new_n698_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n645_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n692_), .A2(new_n334_), .A3(new_n740_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(new_n212_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(new_n645_), .ZN(G1336gat));
  OAI21_X1  g564(.A(new_n202_), .B1(new_n760_), .B2(new_n539_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT111), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n657_), .A2(new_n203_), .A3(new_n205_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n763_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1337gat));
  NOR2_X1   g569(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n771_));
  OAI21_X1  g570(.A(G99gat), .B1(new_n763_), .B2(new_n594_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n761_), .A2(new_n222_), .A3(new_n558_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n774_), .B(new_n775_), .Z(G1338gat));
  OAI21_X1  g575(.A(G106gat), .B1(new_n763_), .B2(new_n449_), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n778_));
  XNOR2_X1  g577(.A(new_n777_), .B(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n761_), .A2(new_n223_), .A3(new_n672_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n612_), .A2(new_n638_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n633_), .B2(new_n787_), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT114), .B(KEYINPUT55), .C1(new_n629_), .C2(new_n632_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n628_), .A2(new_n787_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n630_), .A2(new_n620_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n622_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n788_), .A2(new_n789_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n617_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n633_), .A2(new_n787_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT114), .ZN(new_n798_));
  INV_X1    g597(.A(new_n793_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n633_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n617_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n785_), .B1(new_n796_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n596_), .A2(new_n601_), .A3(new_n598_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n600_), .A2(new_n597_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n605_), .A3(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n609_), .B(new_n807_), .C1(new_n640_), .C2(new_n636_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n648_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n783_), .B1(new_n809_), .B2(KEYINPUT57), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n795_), .B1(new_n794_), .B2(new_n617_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n802_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n784_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n808_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT57), .B(new_n299_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n609_), .A2(new_n638_), .A3(new_n807_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n796_), .B2(new_n803_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI221_X1 g620(.A(new_n818_), .B1(KEYINPUT117), .B2(KEYINPUT58), .C1(new_n796_), .C2(new_n803_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n684_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n299_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(KEYINPUT115), .A3(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n810_), .A2(new_n815_), .A3(new_n823_), .A4(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n612_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n303_), .A2(new_n828_), .A3(new_n739_), .A4(new_n335_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT54), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n829_), .A2(KEYINPUT54), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n827_), .A2(new_n334_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n672_), .A2(new_n657_), .A3(new_n594_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n645_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n612_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n824_), .A2(new_n825_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n823_), .A2(new_n837_), .A3(new_n815_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n334_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n831_), .A2(new_n830_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n834_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n842_), .A2(KEYINPUT118), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT59), .B1(new_n842_), .B2(KEYINPUT118), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT119), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n841_), .A2(new_n847_), .A3(new_n843_), .A4(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n832_), .B2(new_n834_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n849_), .A2(new_n828_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n836_), .B1(new_n852_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g652(.A(new_n739_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n846_), .A2(new_n854_), .A3(new_n850_), .A4(new_n848_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G120gat), .ZN(new_n856_));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n739_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n835_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n857_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n856_), .A2(KEYINPUT120), .A3(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1341gat));
  AOI21_X1  g663(.A(G127gat), .B1(new_n835_), .B2(new_n335_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n849_), .A2(new_n342_), .A3(new_n851_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n335_), .ZN(G1342gat));
  INV_X1    g666(.A(new_n835_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n343_), .B1(new_n868_), .B2(new_n299_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n846_), .A2(G134gat), .A3(new_n850_), .A4(new_n848_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n303_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT121), .ZN(G1343gat));
  NOR2_X1   g671(.A1(new_n832_), .A2(new_n657_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n449_), .A2(new_n558_), .A3(new_n404_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n828_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n360_), .ZN(G1344gat));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n739_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n361_), .ZN(G1345gat));
  NOR2_X1   g678(.A1(new_n875_), .A2(new_n334_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT61), .B(G155gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  NOR3_X1   g681(.A1(new_n875_), .A2(new_n282_), .A3(new_n303_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n873_), .A2(new_n648_), .A3(new_n874_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n282_), .B2(new_n884_), .ZN(G1347gat));
  NOR3_X1   g684(.A1(new_n594_), .A2(new_n539_), .A3(new_n645_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n886_), .A2(new_n449_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n841_), .A2(new_n612_), .A3(new_n887_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n888_), .A2(G169gat), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n889_), .A2(KEYINPUT122), .A3(new_n890_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n893_), .B(new_n894_), .C1(new_n890_), .C2(new_n889_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n841_), .A2(new_n887_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT123), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n612_), .B1(new_n475_), .B2(new_n474_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n895_), .B1(new_n897_), .B2(new_n898_), .ZN(G1348gat));
  INV_X1    g698(.A(new_n897_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G176gat), .B1(new_n900_), .B2(new_n854_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n832_), .A2(new_n672_), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n854_), .A2(new_n886_), .A3(G176gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1349gat));
  NOR3_X1   g703(.A1(new_n897_), .A2(new_n469_), .A3(new_n334_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n902_), .A2(new_n335_), .A3(new_n886_), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT124), .Z(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n907_), .B2(new_n482_), .ZN(G1350gat));
  OAI21_X1  g707(.A(G190gat), .B1(new_n897_), .B2(new_n303_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n648_), .A2(new_n468_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n897_), .B2(new_n910_), .ZN(G1351gat));
  NAND2_X1  g710(.A1(new_n594_), .A2(new_n590_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(KEYINPUT125), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n832_), .A2(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n539_), .B1(new_n912_), .B2(KEYINPUT125), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n828_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(new_n420_), .ZN(G1352gat));
  INV_X1    g717(.A(new_n916_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n854_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n412_), .A2(KEYINPUT126), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1353gat));
  NOR2_X1   g721(.A1(new_n916_), .A2(new_n334_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n923_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924_));
  XOR2_X1   g723(.A(KEYINPUT63), .B(G211gat), .Z(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n923_), .B2(new_n925_), .ZN(G1354gat));
  NAND3_X1  g725(.A1(new_n919_), .A2(KEYINPUT127), .A3(new_n648_), .ZN(new_n927_));
  INV_X1    g726(.A(G218gat), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(new_n916_), .B2(new_n299_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n928_), .A3(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n919_), .A2(G218gat), .A3(new_n684_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1355gat));
endmodule


