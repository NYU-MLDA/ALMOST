//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n805_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_;
  AND2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n205_), .A2(KEYINPUT84), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT79), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G183gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n208_), .B1(new_n213_), .B2(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n205_), .A2(KEYINPUT84), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n206_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT83), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT25), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT80), .B1(new_n222_), .B2(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n224_));
  INV_X1    g023(.A(G190gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT26), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT81), .B1(new_n225_), .B2(KEYINPUT26), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT81), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(new_n222_), .A3(G190gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n221_), .A2(new_n227_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT82), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n221_), .A2(new_n234_), .A3(new_n231_), .A4(new_n227_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n202_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n218_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  AOI211_X1 g040(.A(KEYINPUT83), .B(new_n239_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n238_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n208_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n217_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G127gat), .B(G134gat), .Z(new_n247_));
  XOR2_X1   g046(.A(G113gat), .B(G120gat), .Z(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  INV_X1    g048(.A(KEYINPUT85), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT85), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT30), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n246_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT31), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n255_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G15gat), .B(G43gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G71gat), .B(G99gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G197gat), .B(G204gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n265_), .A2(KEYINPUT21), .B1(new_n266_), .B2(KEYINPUT87), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n265_), .B2(KEYINPUT21), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270_));
  OR2_X1    g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n272_), .B(KEYINPUT3), .Z(new_n273_));
  NAND2_X1  g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT2), .Z(new_n275_));
  OAI211_X1 g074(.A(new_n270_), .B(new_n271_), .C1(new_n273_), .C2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n272_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n270_), .A2(KEYINPUT1), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n271_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n270_), .A2(KEYINPUT1), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n277_), .B(new_n274_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n269_), .B1(KEYINPUT29), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G228gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G78gat), .B(G106gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT88), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n282_), .A2(KEYINPUT29), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G22gat), .B(G50gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n285_), .A2(new_n286_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT89), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(KEYINPUT89), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n288_), .A2(new_n293_), .A3(new_n295_), .A4(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n287_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(new_n294_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(new_n293_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G8gat), .B(G36gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G92gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT18), .B(G64gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n205_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT90), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n222_), .A2(G190gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n225_), .A2(KEYINPUT26), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT25), .B(G183gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n245_), .A2(new_n240_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n269_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT20), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT19), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT91), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n228_), .A2(new_n230_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n220_), .B2(new_n219_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n234_), .B1(new_n325_), .B2(new_n227_), .ZN(new_n326_));
  AND4_X1   g125(.A1(new_n234_), .A2(new_n221_), .A3(new_n227_), .A4(new_n231_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n240_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT83), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n236_), .A2(new_n218_), .A3(new_n240_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n245_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n216_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n323_), .B1(new_n332_), .B2(new_n318_), .ZN(new_n333_));
  AOI211_X1 g132(.A(KEYINPUT91), .B(new_n269_), .C1(new_n331_), .C2(new_n216_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n322_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n321_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n331_), .A2(new_n216_), .A3(new_n269_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT20), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n307_), .B1(new_n335_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n335_), .A2(new_n341_), .A3(new_n307_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT92), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT92), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n342_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n253_), .A2(new_n282_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT93), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT4), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n282_), .A2(new_n249_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n253_), .B2(new_n282_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT4), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n350_), .B1(new_n349_), .B2(KEYINPUT4), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n351_), .A2(new_n353_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G85gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT0), .B(G57gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  NAND2_X1  g161(.A1(new_n355_), .A2(new_n352_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT94), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(KEYINPUT33), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n351_), .A2(new_n352_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n362_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n355_), .A2(new_n353_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n371_), .A2(KEYINPUT95), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n364_), .A2(new_n366_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(KEYINPUT95), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n367_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n345_), .A2(new_n348_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n358_), .A2(new_n363_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n369_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n364_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT91), .B1(new_n246_), .B2(new_n269_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n332_), .A2(new_n323_), .A3(new_n318_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n383_));
  AND2_X1   g182(.A1(new_n269_), .A2(new_n316_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(new_n309_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n336_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n337_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT97), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n307_), .A2(KEYINPUT32), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n379_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n340_), .B1(new_n382_), .B2(new_n322_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n391_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n302_), .B1(new_n376_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT98), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n387_), .B(KEYINPUT97), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n385_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n321_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n307_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n344_), .A2(KEYINPUT27), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n396_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n306_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT27), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n393_), .B2(new_n307_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n405_), .A3(KEYINPUT98), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n379_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT27), .B1(new_n343_), .B2(new_n344_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n407_), .A2(new_n408_), .A3(new_n301_), .A4(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n264_), .B1(new_n395_), .B2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT98), .B1(new_n403_), .B2(new_n405_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n400_), .A2(new_n401_), .A3(new_n396_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n410_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n407_), .A2(KEYINPUT99), .A3(new_n410_), .ZN(new_n418_));
  AOI211_X1 g217(.A(new_n379_), .B(new_n301_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT100), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT100), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n417_), .A2(new_n418_), .A3(new_n422_), .A4(new_n419_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n412_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G1gat), .B(G8gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT76), .Z(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT75), .B(G1gat), .ZN(new_n427_));
  INV_X1    g226(.A(G8gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT14), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G15gat), .B(G22gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n426_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G29gat), .B(G36gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G43gat), .B(G50gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n432_), .B(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(G229gat), .A3(G233gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n435_), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n435_), .B(KEYINPUT15), .Z(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n432_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G229gat), .A2(G233gat), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT77), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n437_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G113gat), .B(G141gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G169gat), .B(G197gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT78), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n444_), .A2(new_n447_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT7), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT6), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G85gat), .B(G92gat), .Z(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT8), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT8), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT65), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n457_), .B(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n464_), .A2(new_n455_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT66), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n462_), .B(new_n459_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n465_), .A2(new_n466_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n461_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT64), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT9), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n459_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT10), .B(G99gat), .Z(new_n475_));
  INV_X1    g274(.A(G106gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n471_), .A2(new_n472_), .A3(G85gat), .A4(G92gat), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n464_), .A2(new_n474_), .A3(new_n477_), .A4(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n469_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G71gat), .B(G78gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(G57gat), .B(G64gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT11), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n482_), .A2(KEYINPUT11), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n481_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n481_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n483_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(KEYINPUT12), .A3(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT68), .Z(new_n491_));
  XOR2_X1   g290(.A(new_n489_), .B(KEYINPUT67), .Z(new_n492_));
  NOR2_X1   g291(.A1(new_n480_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n492_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n469_), .B2(new_n479_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n495_), .A2(KEYINPUT70), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT70), .B1(new_n495_), .B2(new_n497_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n493_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G230gat), .A2(G233gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n491_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(G230gat), .B(G233gat), .C1(new_n493_), .C2(new_n495_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT5), .B(G176gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(G204gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G120gat), .B(G148gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n502_), .A2(new_n503_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT13), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n512_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n424_), .A2(new_n453_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G231gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n432_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(new_n492_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G127gat), .B(G155gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G211gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT16), .B(G183gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n523_), .B(KEYINPUT17), .Z(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n518_), .A2(new_n489_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n518_), .A2(new_n489_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n526_), .A2(KEYINPUT17), .A3(new_n523_), .A4(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n533_), .A2(KEYINPUT35), .ZN(new_n534_));
  INV_X1    g333(.A(new_n480_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n535_), .A2(KEYINPUT72), .A3(new_n435_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT72), .B1(new_n535_), .B2(new_n435_), .ZN(new_n537_));
  OAI221_X1 g336(.A(new_n534_), .B1(new_n439_), .B2(new_n535_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n533_), .A2(KEYINPUT35), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G190gat), .B(G218gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT36), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT74), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n544_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT73), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n540_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT37), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n516_), .A2(new_n530_), .A3(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n379_), .A3(new_n427_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT101), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT38), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n547_), .A2(KEYINPUT102), .A3(new_n550_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT102), .B1(new_n547_), .B2(new_n550_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n516_), .A2(new_n530_), .A3(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(G1gat), .B1(new_n564_), .B2(new_n408_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n565_), .ZN(G1324gat));
  AOI21_X1  g365(.A(KEYINPUT99), .B1(new_n407_), .B2(new_n410_), .ZN(new_n567_));
  AOI211_X1 g366(.A(new_n416_), .B(new_n409_), .C1(new_n402_), .C2(new_n406_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(G8gat), .B1(new_n564_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT39), .ZN(new_n571_));
  INV_X1    g370(.A(new_n569_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n556_), .A2(new_n428_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(G1325gat));
  INV_X1    g375(.A(new_n264_), .ZN(new_n577_));
  OAI21_X1  g376(.A(G15gat), .B1(new_n564_), .B2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT41), .Z(new_n579_));
  INV_X1    g378(.A(G15gat), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n556_), .A2(new_n580_), .A3(new_n264_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(G1326gat));
  OAI21_X1  g381(.A(G22gat), .B1(new_n564_), .B2(new_n302_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT42), .ZN(new_n584_));
  INV_X1    g383(.A(G22gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n556_), .A2(new_n585_), .A3(new_n301_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT104), .ZN(G1327gat));
  NOR2_X1   g387(.A1(new_n563_), .A2(new_n530_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n516_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(G29gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n379_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n412_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n422_), .B1(new_n569_), .B2(new_n419_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n423_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n555_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n594_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT105), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT43), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n424_), .A2(new_n555_), .A3(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n515_), .A2(new_n453_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n604_), .A2(KEYINPUT44), .A3(new_n605_), .A4(new_n529_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n598_), .A2(new_n601_), .A3(new_n599_), .A4(KEYINPUT43), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n593_), .B1(new_n424_), .B2(new_n555_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n605_), .A4(new_n529_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT44), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(new_n379_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n592_), .B1(new_n613_), .B2(new_n591_), .ZN(G1328gat));
  NAND3_X1  g413(.A1(new_n606_), .A2(new_n572_), .A3(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT106), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT106), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n606_), .A2(new_n617_), .A3(new_n611_), .A4(new_n572_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(G36gat), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT107), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT107), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n616_), .A2(new_n621_), .A3(G36gat), .A4(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(G36gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n590_), .A2(new_n624_), .A3(new_n572_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT108), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT45), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n623_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n623_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1329gat));
  NAND2_X1  g432(.A1(new_n612_), .A2(new_n264_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n577_), .A2(G43gat), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n634_), .A2(G43gat), .B1(new_n590_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g436(.A(G50gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n590_), .A2(new_n638_), .A3(new_n301_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT110), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n612_), .A2(new_n301_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(G50gat), .ZN(new_n642_));
  AOI211_X1 g441(.A(KEYINPUT110), .B(new_n638_), .C1(new_n612_), .C2(new_n301_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(G1331gat));
  AND2_X1   g443(.A1(new_n513_), .A2(new_n514_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n452_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n424_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n530_), .A3(new_n555_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT111), .ZN(new_n650_));
  AOI21_X1  g449(.A(G57gat), .B1(new_n650_), .B2(new_n379_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n530_), .A3(new_n563_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n408_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(G57gat), .B2(new_n653_), .ZN(G1332gat));
  OAI21_X1  g453(.A(G64gat), .B1(new_n652_), .B2(new_n569_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT48), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n569_), .A2(G64gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT112), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n650_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n659_), .ZN(G1333gat));
  OAI21_X1  g459(.A(G71gat), .B1(new_n652_), .B2(new_n577_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT49), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n577_), .A2(G71gat), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT113), .Z(new_n664_));
  NAND2_X1  g463(.A1(new_n650_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(G1334gat));
  OAI21_X1  g465(.A(G78gat), .B1(new_n652_), .B2(new_n302_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT50), .ZN(new_n668_));
  INV_X1    g467(.A(G78gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n650_), .A2(new_n669_), .A3(new_n301_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1335gat));
  NAND2_X1  g470(.A1(new_n648_), .A2(new_n589_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT114), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G85gat), .B1(new_n674_), .B2(new_n379_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n604_), .A2(KEYINPUT115), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n604_), .A2(KEYINPUT115), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(new_n529_), .A3(new_n646_), .A4(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n408_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n675_), .B1(new_n679_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g479(.A(G92gat), .B1(new_n674_), .B2(new_n572_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n678_), .A2(new_n569_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g482(.A(G99gat), .B1(new_n678_), .B2(new_n577_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n674_), .A2(new_n475_), .A3(new_n264_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n686_), .B(new_n687_), .Z(G1338gat));
  NAND3_X1  g487(.A1(new_n604_), .A2(new_n301_), .A3(new_n529_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G106gat), .B1(new_n689_), .B2(new_n647_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n690_), .A2(KEYINPUT52), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(KEYINPUT52), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n302_), .A2(G106gat), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n691_), .A2(new_n692_), .B1(new_n674_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n694_), .B(new_n695_), .Z(G1339gat));
  NOR2_X1   g495(.A1(new_n577_), .A2(new_n301_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n572_), .A2(new_n408_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n501_), .B1(new_n491_), .B2(new_n500_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT55), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n502_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n491_), .A2(new_n500_), .A3(KEYINPUT55), .A4(new_n501_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(KEYINPUT56), .A3(new_n507_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT120), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n508_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n703_), .A2(new_n507_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT56), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n706_), .A2(new_n708_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n509_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n452_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n436_), .A2(new_n442_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(new_n447_), .C1(new_n440_), .C2(new_n442_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n448_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n511_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT121), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n714_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT57), .B1(new_n721_), .B2(new_n563_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT57), .ZN(new_n723_));
  AOI211_X1 g522(.A(new_n723_), .B(new_n562_), .C1(new_n714_), .C2(new_n720_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n704_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n707_), .A2(KEYINPUT56), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n713_), .B(new_n717_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT58), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n599_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n530_), .B1(new_n725_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT119), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n452_), .A2(new_n529_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n645_), .B1(KEYINPUT118), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(KEYINPUT118), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n555_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n732_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT118), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n515_), .B1(new_n739_), .B2(new_n733_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n740_), .A2(KEYINPUT119), .A3(new_n555_), .A4(new_n736_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n741_), .A3(KEYINPUT54), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT54), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n732_), .B(new_n743_), .C1(new_n735_), .C2(new_n737_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n697_), .B(new_n698_), .C1(new_n731_), .C2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G113gat), .B1(new_n747_), .B2(new_n452_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n721_), .A2(new_n563_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n723_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n721_), .A2(KEYINPUT57), .A3(new_n563_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n730_), .A3(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n529_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n742_), .A2(new_n744_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n758_));
  NAND4_X1  g557(.A1(new_n757_), .A2(new_n697_), .A3(new_n698_), .A4(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n750_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(G113gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n748_), .B1(new_n761_), .B2(new_n452_), .ZN(G1340gat));
  INV_X1    g561(.A(G120gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n645_), .B2(KEYINPUT60), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n747_), .B(new_n764_), .C1(KEYINPUT60), .C2(new_n763_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n645_), .B1(new_n750_), .B2(new_n759_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n763_), .ZN(G1341gat));
  AOI21_X1  g566(.A(G127gat), .B1(new_n747_), .B2(new_n530_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n530_), .A2(G127gat), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT123), .Z(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n760_), .B2(new_n770_), .ZN(G1342gat));
  INV_X1    g570(.A(KEYINPUT124), .ZN(new_n772_));
  INV_X1    g571(.A(G134gat), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n773_), .B(new_n555_), .C1(new_n750_), .C2(new_n759_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G134gat), .B1(new_n747_), .B2(new_n562_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n772_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n760_), .A2(G134gat), .A3(new_n599_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n775_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(KEYINPUT124), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(G1343gat));
  AOI211_X1 g579(.A(new_n264_), .B(new_n302_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n698_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(new_n453_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g583(.A1(new_n782_), .A2(new_n645_), .ZN(new_n785_));
  XOR2_X1   g584(.A(KEYINPUT125), .B(G148gat), .Z(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(G1345gat));
  NOR2_X1   g586(.A1(new_n782_), .A2(new_n529_), .ZN(new_n788_));
  XOR2_X1   g587(.A(KEYINPUT61), .B(G155gat), .Z(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(G1346gat));
  INV_X1    g589(.A(G162gat), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n782_), .A2(new_n791_), .A3(new_n555_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n781_), .A2(new_n562_), .A3(new_n698_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n791_), .B2(new_n793_), .ZN(G1347gat));
  NOR2_X1   g593(.A1(new_n569_), .A2(new_n379_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n757_), .A2(new_n697_), .A3(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G169gat), .B1(new_n796_), .B2(new_n453_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(KEYINPUT62), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(KEYINPUT62), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n452_), .A2(new_n203_), .ZN(new_n800_));
  XOR2_X1   g599(.A(new_n800_), .B(KEYINPUT126), .Z(new_n801_));
  OAI22_X1  g600(.A1(new_n798_), .A2(new_n799_), .B1(new_n796_), .B2(new_n801_), .ZN(G1348gat));
  NOR2_X1   g601(.A1(new_n796_), .A2(new_n645_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(new_n204_), .ZN(G1349gat));
  NOR2_X1   g603(.A1(new_n796_), .A2(new_n529_), .ZN(new_n805_));
  MUX2_X1   g604(.A(new_n213_), .B(new_n314_), .S(new_n805_), .Z(G1350gat));
  OAI21_X1  g605(.A(G190gat), .B1(new_n796_), .B2(new_n555_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n757_), .A2(new_n313_), .A3(new_n697_), .A4(new_n795_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n563_), .B2(new_n808_), .ZN(G1351gat));
  NAND2_X1  g608(.A1(new_n781_), .A2(new_n795_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n453_), .ZN(new_n811_));
  XOR2_X1   g610(.A(new_n811_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n645_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(G204gat), .Z(G1353gat));
  NAND3_X1  g613(.A1(new_n781_), .A2(new_n530_), .A3(new_n795_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n816_));
  AND2_X1   g615(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n815_), .B2(new_n816_), .ZN(G1354gat));
  INV_X1    g618(.A(G218gat), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n810_), .A2(new_n820_), .A3(new_n555_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n781_), .A2(new_n562_), .A3(new_n795_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(new_n822_), .ZN(G1355gat));
endmodule


