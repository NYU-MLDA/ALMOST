//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_, new_n954_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT69), .ZN(new_n203_));
  XOR2_X1   g002(.A(G43gat), .B(G50gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT15), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT10), .B(G99gat), .Z(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(KEYINPUT64), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n214_), .B(new_n215_), .C1(KEYINPUT64), .C2(KEYINPUT9), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n218_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n210_), .A2(new_n213_), .A3(new_n216_), .A4(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n212_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n208_), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n222_), .B(new_n225_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n215_), .A2(new_n217_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT8), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n228_), .A2(new_n231_), .A3(new_n229_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n218_), .A2(new_n230_), .A3(new_n219_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n228_), .A2(new_n229_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n221_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n206_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT35), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G232gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT34), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n238_), .A2(new_n205_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(new_n239_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G190gat), .B(G218gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(G134gat), .B(G162gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT71), .Z(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n251_), .B(KEYINPUT36), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT37), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n255_), .A2(KEYINPUT37), .A3(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G127gat), .B(G155gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT16), .ZN(new_n266_));
  XOR2_X1   g065(.A(G183gat), .B(G211gat), .Z(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(KEYINPUT17), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT17), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT73), .B(G1gat), .ZN(new_n272_));
  INV_X1    g071(.A(G8gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT14), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT72), .B(G15gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(G22gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G1gat), .B(G8gat), .Z(new_n280_));
  OR2_X1    g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G231gat), .A2(G233gat), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n283_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G71gat), .B(G78gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(G57gat), .B(G64gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n286_), .B1(KEYINPUT11), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n287_), .B2(KEYINPUT11), .ZN(new_n290_));
  INV_X1    g089(.A(G64gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G57gat), .ZN(new_n292_));
  INV_X1    g091(.A(G57gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G64gat), .ZN(new_n294_));
  AND4_X1   g093(.A1(new_n289_), .A2(new_n292_), .A3(new_n294_), .A4(KEYINPUT11), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n288_), .B1(new_n290_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n294_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT11), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT66), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n287_), .A2(new_n289_), .A3(KEYINPUT11), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n298_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .A4(new_n286_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n284_), .A2(new_n285_), .A3(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n296_), .A2(new_n302_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n282_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n279_), .A2(new_n280_), .ZN(new_n307_));
  OAI211_X1 g106(.A(G231gat), .B(G233gat), .C1(new_n306_), .C2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n305_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n271_), .B1(new_n304_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n270_), .B1(new_n311_), .B2(new_n269_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n303_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n308_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n312_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n316_), .B1(new_n304_), .B2(new_n310_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT76), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n268_), .B1(new_n315_), .B2(new_n271_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n323_), .B(new_n318_), .C1(new_n324_), .C2(new_n270_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n264_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT77), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n281_), .A2(new_n282_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(new_n205_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G229gat), .A2(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n206_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n205_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n331_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G113gat), .B(G141gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(G169gat), .B(G197gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n333_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT12), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n236_), .A2(new_n305_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n225_), .A2(new_n222_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n229_), .B1(new_n209_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n231_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n228_), .A2(new_n231_), .A3(new_n229_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n303_), .A3(new_n221_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n344_), .B1(new_n345_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G230gat), .A2(G233gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT12), .B1(new_n236_), .B2(new_n305_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n353_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n345_), .B2(new_n352_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G176gat), .B(G204gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT68), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G120gat), .B(G148gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n357_), .A2(new_n358_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT13), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(KEYINPUT13), .A3(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n343_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT25), .B(G183gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT78), .B(G190gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT26), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT23), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT24), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  MUX2_X1   g184(.A(new_n384_), .B(KEYINPUT24), .S(new_n385_), .Z(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n382_), .A3(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT80), .B(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT22), .ZN(new_n389_));
  OAI21_X1  g188(.A(G169gat), .B1(new_n389_), .B2(KEYINPUT79), .ZN(new_n390_));
  INV_X1    g189(.A(G169gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT22), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n388_), .B(new_n390_), .C1(KEYINPUT79), .C2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(G183gat), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n376_), .A2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n381_), .B(KEYINPUT23), .Z(new_n396_));
  OAI211_X1 g195(.A(new_n393_), .B(new_n383_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n387_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G71gat), .B(G99gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G43gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n398_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(G15gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT30), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n401_), .B(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n406_), .A2(KEYINPUT82), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(KEYINPUT82), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G113gat), .B(G120gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G127gat), .B(G134gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT81), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n411_), .A2(KEYINPUT81), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n410_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n411_), .A2(KEYINPUT81), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT31), .ZN(new_n419_));
  OR3_X1    g218(.A1(new_n407_), .A2(new_n408_), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n406_), .A2(KEYINPUT82), .A3(new_n419_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT18), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G64gat), .B(G92gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n424_), .B(new_n425_), .Z(new_n426_));
  XNOR2_X1  g225(.A(G197gat), .B(G204gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G211gat), .B(G218gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n428_), .B(KEYINPUT86), .Z(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT21), .B(new_n427_), .C1(new_n429_), .C2(KEYINPUT87), .ZN(new_n430_));
  INV_X1    g229(.A(new_n427_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n429_), .B2(KEYINPUT21), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT21), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n428_), .B(KEYINPUT86), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n430_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n398_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT19), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT22), .B(G169gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n388_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n443_), .B(new_n383_), .C1(new_n396_), .C2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT26), .B(G190gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n375_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n386_), .A2(new_n382_), .A3(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n430_), .B(new_n449_), .C1(new_n432_), .C2(new_n436_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n438_), .A2(KEYINPUT20), .A3(new_n441_), .A4(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n452_));
  INV_X1    g251(.A(new_n449_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n452_), .B1(new_n437_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n398_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n455_), .B(new_n430_), .C1(new_n436_), .C2(new_n432_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n440_), .B(KEYINPUT90), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n426_), .B(new_n451_), .C1(new_n457_), .C2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT27), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n454_), .A2(new_n459_), .A3(new_n456_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n450_), .A2(KEYINPUT20), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n450_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n438_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n462_), .B1(new_n467_), .B2(new_n440_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT96), .B1(new_n468_), .B2(new_n426_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT96), .ZN(new_n470_));
  INV_X1    g269(.A(new_n426_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n463_), .A2(new_n464_), .B1(new_n437_), .B2(new_n398_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n441_), .B1(new_n472_), .B2(new_n466_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n470_), .B(new_n471_), .C1(new_n473_), .C2(new_n462_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n461_), .B1(new_n469_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n451_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n459_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n471_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT27), .B1(new_n460_), .B2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G1gat), .B(G29gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G85gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  NOR2_X1   g284(.A1(G155gat), .A2(G162gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G155gat), .A2(G162gat), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n486_), .B1(new_n491_), .B2(KEYINPUT1), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT1), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n493_), .A3(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G141gat), .A2(G148gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(G141gat), .A2(G148gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n498_), .B(KEYINPUT3), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n496_), .B(KEYINPUT2), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n486_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT4), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n418_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G225gat), .A2(G233gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n418_), .A2(new_n506_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n495_), .A2(new_n499_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n415_), .A2(new_n417_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT91), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n418_), .A2(new_n506_), .A3(KEYINPUT91), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT4), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(KEYINPUT92), .A3(KEYINPUT4), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n511_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n509_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n485_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT92), .B1(new_n518_), .B2(KEYINPUT4), .ZN(new_n528_));
  AOI211_X1 g327(.A(new_n520_), .B(new_n507_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n510_), .B(new_n508_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n485_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n524_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n526_), .A2(new_n527_), .A3(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n530_), .A2(KEYINPUT95), .A3(new_n524_), .A4(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G78gat), .B(G106gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n506_), .A2(KEYINPUT29), .ZN(new_n537_));
  INV_X1    g336(.A(G233gat), .ZN(new_n538_));
  NOR2_X1   g337(.A1(KEYINPUT85), .A2(G228gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(KEYINPUT85), .A2(G228gat), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n437_), .A2(new_n537_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n437_), .B2(new_n537_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n536_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n437_), .A2(new_n537_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n542_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n536_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n544_), .A3(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n551_), .A3(KEYINPUT88), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT84), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT28), .B1(new_n506_), .B2(KEYINPUT29), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT28), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT29), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n513_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n553_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G22gat), .B(G50gat), .Z(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n553_), .A3(new_n557_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n560_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n561_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n563_), .B1(new_n564_), .B2(new_n558_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT88), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n549_), .A2(new_n566_), .A3(new_n544_), .A4(new_n550_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n552_), .A2(new_n562_), .A3(new_n565_), .A4(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n562_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT89), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n547_), .A2(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT89), .B(new_n536_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n569_), .A2(new_n571_), .A3(new_n572_), .A4(new_n551_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n480_), .A2(new_n535_), .A3(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n426_), .A2(KEYINPUT32), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n476_), .A2(new_n477_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n468_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n579_), .B2(new_n577_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n533_), .A2(new_n534_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n460_), .A2(new_n478_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n509_), .B(new_n508_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n531_), .B1(new_n518_), .B2(new_n510_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT33), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n532_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n530_), .A2(KEYINPUT33), .A3(new_n524_), .A4(new_n531_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n575_), .B1(new_n581_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n422_), .B1(new_n576_), .B2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n533_), .A2(new_n534_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n422_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n574_), .A3(new_n480_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n374_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n328_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n592_), .A3(new_n272_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT38), .ZN(new_n598_));
  INV_X1    g397(.A(new_n259_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n321_), .A2(new_n325_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n374_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n592_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(G1gat), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n598_), .A2(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(new_n480_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n596_), .A2(new_n273_), .A3(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n610_), .B(new_n606_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n612_), .A2(new_n613_), .A3(G8gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n612_), .B2(G8gat), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(G1325gat));
  INV_X1    g417(.A(new_n422_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n604_), .A2(new_n619_), .A3(new_n606_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G15gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n596_), .A2(new_n403_), .A3(new_n619_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(G1326gat));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n596_), .A2(new_n627_), .A3(new_n575_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n604_), .A2(new_n575_), .A3(new_n606_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT42), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(new_n630_), .A3(G22gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n629_), .B2(G22gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(G1327gat));
  NOR2_X1   g432(.A1(new_n326_), .A2(new_n259_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n595_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n592_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n263_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n581_), .A2(new_n589_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n475_), .A2(new_n574_), .A3(new_n479_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n642_), .A2(new_n574_), .B1(new_n643_), .B2(new_n535_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n594_), .B1(new_n644_), .B2(new_n619_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n264_), .A2(KEYINPUT99), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n263_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n645_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n641_), .B1(new_n650_), .B2(KEYINPUT43), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n605_), .A2(new_n373_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n638_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n640_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n645_), .A2(new_n654_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n591_), .A2(new_n594_), .B1(new_n648_), .B2(new_n646_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(new_n639_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n657_), .A2(KEYINPUT44), .A3(new_n373_), .A4(new_n605_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n653_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n592_), .A2(G29gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n637_), .B1(new_n659_), .B2(new_n660_), .ZN(G1328gat));
  NOR2_X1   g460(.A1(new_n480_), .A2(G36gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n595_), .A2(new_n634_), .A3(new_n662_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(KEYINPUT100), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(KEYINPUT100), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(KEYINPUT45), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT45), .B1(new_n664_), .B2(new_n665_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n653_), .A2(new_n658_), .A3(new_n610_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G36gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n668_), .A2(KEYINPUT46), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1329gat));
  NAND4_X1  g474(.A1(new_n653_), .A2(new_n658_), .A3(G43gat), .A4(new_n619_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT101), .B(G43gat), .Z(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(new_n635_), .B2(new_n422_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g479(.A(G50gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n636_), .A2(new_n681_), .A3(new_n575_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n659_), .A2(new_n575_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(G50gat), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT102), .B(new_n681_), .C1(new_n659_), .C2(new_n575_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(G1331gat));
  NAND2_X1  g486(.A1(new_n343_), .A2(new_n372_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n328_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n592_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT103), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n605_), .A2(new_n688_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n604_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n535_), .A2(new_n293_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n692_), .B1(new_n694_), .B2(new_n695_), .ZN(G1332gat));
  NAND3_X1  g495(.A1(new_n690_), .A2(new_n291_), .A3(new_n610_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n610_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(G64gat), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT48), .B(new_n291_), .C1(new_n694_), .C2(new_n610_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1333gat));
  INV_X1    g501(.A(G71gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n690_), .A2(new_n703_), .A3(new_n619_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n694_), .A2(new_n619_), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(G71gat), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G71gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(G1334gat));
  INV_X1    g508(.A(G78gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n690_), .A2(new_n710_), .A3(new_n575_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n694_), .A2(new_n575_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(G78gat), .ZN(new_n714_));
  AOI211_X1 g513(.A(KEYINPUT50), .B(new_n710_), .C1(new_n694_), .C2(new_n575_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(G1335gat));
  NAND2_X1  g515(.A1(new_n689_), .A2(new_n634_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n689_), .A2(KEYINPUT105), .A3(new_n634_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G85gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n592_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n657_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n688_), .A2(new_n326_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n655_), .B(KEYINPUT106), .C1(new_n656_), .C2(new_n639_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n592_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n723_), .B1(new_n729_), .B2(new_n722_), .ZN(G1336gat));
  INV_X1    g529(.A(G92gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n721_), .A2(new_n731_), .A3(new_n610_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n728_), .A2(new_n610_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n731_), .ZN(G1337gat));
  NAND4_X1  g533(.A1(new_n725_), .A2(new_n727_), .A3(new_n619_), .A4(new_n726_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n619_), .A2(new_n211_), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n735_), .A2(G99gat), .B1(new_n721_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT107), .ZN(new_n740_));
  NAND2_X1  g539(.A1(KEYINPUT107), .A2(KEYINPUT51), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743_));
  AOI22_X1  g542(.A1(new_n740_), .A2(new_n742_), .B1(new_n743_), .B2(new_n739_), .ZN(G1338gat));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n721_), .A2(new_n212_), .A3(new_n575_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT110), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n688_), .A2(new_n326_), .A3(new_n574_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n639_), .B1(new_n645_), .B2(new_n649_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT109), .B(new_n750_), .C1(new_n751_), .C2(new_n641_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G106gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT109), .B1(new_n657_), .B2(new_n750_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n749_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756_));
  INV_X1    g555(.A(new_n750_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n651_), .B2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n758_), .A2(G106gat), .A3(new_n748_), .A4(new_n752_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n755_), .A2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n747_), .A2(KEYINPUT110), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n745_), .B(new_n746_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n755_), .B2(new_n759_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n746_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT53), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1339gat));
  AOI21_X1  g565(.A(new_n339_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n334_), .A2(new_n335_), .A3(new_n332_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(new_n340_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n366_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n236_), .A2(new_n305_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n303_), .B1(new_n351_), .B2(new_n221_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT12), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n356_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n355_), .A2(KEYINPUT113), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n355_), .A2(KEYINPUT55), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n353_), .A2(new_n356_), .A3(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n780_), .B2(new_n777_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n775_), .A2(new_n354_), .A3(new_n776_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n782_), .A2(KEYINPUT112), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT112), .B1(new_n782_), .B2(new_n783_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n772_), .B(new_n781_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n357_), .B2(KEYINPUT55), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n782_), .A2(KEYINPUT112), .A3(new_n783_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n772_), .B1(new_n791_), .B2(new_n781_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n364_), .B1(new_n787_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT114), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n786_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n364_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n771_), .B1(new_n795_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n263_), .B1(new_n800_), .B2(KEYINPUT58), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n770_), .A2(new_n366_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n364_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n364_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n794_), .B(new_n804_), .C1(new_n797_), .C2(new_n786_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n802_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT116), .B1(new_n801_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n807_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n800_), .A2(KEYINPUT58), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .A4(new_n263_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n366_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n795_), .B2(new_n799_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n770_), .A2(new_n368_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n259_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n809_), .A2(new_n813_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n814_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n816_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT57), .A3(new_n259_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT57), .B1(new_n825_), .B2(new_n259_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n819_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n605_), .B1(new_n822_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n343_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n605_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n372_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n326_), .A2(KEYINPUT111), .A3(new_n834_), .A4(new_n343_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n830_), .B1(new_n836_), .B2(new_n264_), .ZN(new_n837_));
  AOI211_X1 g636(.A(KEYINPUT54), .B(new_n263_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n829_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n610_), .A2(new_n575_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n592_), .A3(new_n619_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n818_), .A2(new_n820_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(new_n826_), .C1(new_n808_), .C2(new_n801_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n605_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n840_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n843_), .A2(KEYINPUT59), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n845_), .A2(KEYINPUT59), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n343_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G113gat), .ZN(new_n854_));
  OR3_X1    g653(.A1(new_n845_), .A2(G113gat), .A3(new_n343_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1340gat));
  AOI211_X1 g655(.A(new_n820_), .B(new_n599_), .C1(new_n824_), .C2(new_n816_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n846_), .B2(KEYINPUT115), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n858_), .A2(new_n813_), .A3(new_n821_), .A4(new_n809_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n839_), .B1(new_n859_), .B2(new_n605_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT59), .B1(new_n860_), .B2(new_n843_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n849_), .A2(new_n850_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n861_), .A2(KEYINPUT117), .A3(new_n372_), .A4(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n843_), .B1(new_n829_), .B2(new_n840_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n372_), .B(new_n862_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n863_), .A2(new_n868_), .A3(G120gat), .ZN(new_n869_));
  INV_X1    g668(.A(G120gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n834_), .B2(KEYINPUT60), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n864_), .B(new_n871_), .C1(KEYINPUT60), .C2(new_n870_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n872_), .ZN(G1341gat));
  INV_X1    g672(.A(G127gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n845_), .B2(new_n605_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT118), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n877_), .B(new_n874_), .C1(new_n845_), .C2(new_n605_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n605_), .A2(new_n874_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n876_), .A2(new_n878_), .B1(new_n851_), .B2(new_n879_), .ZN(G1342gat));
  AOI21_X1  g679(.A(G134gat), .B1(new_n864_), .B2(new_n599_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n881_), .A2(KEYINPUT119), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(KEYINPUT119), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n263_), .A2(G134gat), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n882_), .A2(new_n883_), .B1(new_n851_), .B2(new_n884_), .ZN(G1343gat));
  AND3_X1   g684(.A1(new_n643_), .A2(new_n592_), .A3(new_n422_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n841_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n343_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT120), .B(G141gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n887_), .A2(new_n834_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT121), .B(G148gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1345gat));
  OAI21_X1  g692(.A(KEYINPUT122), .B1(new_n887_), .B2(new_n605_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n841_), .A2(new_n895_), .A3(new_n326_), .A4(new_n886_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n894_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n894_), .B2(new_n896_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1346gat));
  AND4_X1   g699(.A1(G162gat), .A2(new_n841_), .A3(new_n649_), .A4(new_n886_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n841_), .A2(new_n599_), .A3(new_n886_), .ZN(new_n902_));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1347gat));
  NOR2_X1   g703(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n839_), .B1(new_n605_), .B2(new_n847_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n593_), .A2(new_n610_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n575_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n906_), .A2(new_n343_), .A3(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n905_), .B1(new_n910_), .B2(new_n391_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n912_));
  NAND2_X1  g711(.A1(new_n849_), .A2(new_n908_), .ZN(new_n913_));
  OAI211_X1 g712(.A(G169gat), .B(new_n912_), .C1(new_n913_), .C2(new_n343_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n442_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n911_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT124), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n911_), .A2(new_n914_), .A3(new_n918_), .A4(new_n915_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1348gat));
  INV_X1    g719(.A(new_n388_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n906_), .A2(new_n909_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n372_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n923_), .A2(KEYINPUT125), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(KEYINPUT125), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n860_), .A2(new_n575_), .ZN(new_n926_));
  INV_X1    g725(.A(G176gat), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n907_), .A2(new_n927_), .A3(new_n834_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n924_), .A2(new_n925_), .B1(new_n926_), .B2(new_n928_), .ZN(G1349gat));
  NOR3_X1   g728(.A1(new_n913_), .A2(new_n375_), .A3(new_n605_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n926_), .A2(new_n610_), .A3(new_n593_), .A4(new_n326_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n394_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n913_), .B2(new_n264_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n922_), .A2(new_n446_), .A3(new_n599_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1351gat));
  NAND3_X1  g734(.A1(new_n535_), .A2(new_n575_), .A3(new_n422_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n610_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n937_), .B2(new_n936_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n841_), .A2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n852_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n372_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g743(.A1(new_n940_), .A2(new_n326_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  AND2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n945_), .A2(new_n946_), .A3(new_n947_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n945_), .A2(new_n946_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1354gat));
  AND3_X1   g749(.A1(new_n940_), .A2(G218gat), .A3(new_n263_), .ZN(new_n951_));
  AND3_X1   g750(.A1(new_n841_), .A2(new_n599_), .A3(new_n939_), .ZN(new_n952_));
  OR2_X1    g751(.A1(new_n952_), .A2(KEYINPUT127), .ZN(new_n953_));
  AOI21_X1  g752(.A(G218gat), .B1(new_n952_), .B2(KEYINPUT127), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n951_), .B1(new_n953_), .B2(new_n954_), .ZN(G1355gat));
endmodule


