//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_, new_n975_, new_n976_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT36), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G29gat), .B(G36gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT73), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT15), .Z(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G85gat), .B(G92gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n217_), .B2(KEYINPUT9), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n224_), .A2(KEYINPUT64), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT64), .B1(new_n224_), .B2(new_n225_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n218_), .B(new_n223_), .C1(new_n228_), .C2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n221_), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT65), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n220_), .A2(new_n222_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G106gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n233_), .A2(new_n235_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n230_), .B1(new_n242_), .B2(new_n217_), .ZN(new_n243_));
  AOI211_X1 g042(.A(KEYINPUT8), .B(new_n216_), .C1(new_n241_), .C2(new_n223_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n229_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT35), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G232gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT34), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n212_), .A2(new_n245_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n246_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n253_), .ZN(new_n254_));
  OAI211_X1 g053(.A(KEYINPUT66), .B(new_n229_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n211_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(new_n252_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n252_), .B1(new_n250_), .B2(new_n257_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n207_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT76), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(KEYINPUT76), .B(new_n207_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n260_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT36), .B1(new_n204_), .B2(new_n205_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n258_), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n261_), .A2(new_n269_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT77), .B(KEYINPUT37), .Z(new_n273_));
  AOI22_X1  g072(.A1(new_n270_), .A2(KEYINPUT37), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G231gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT78), .B(G8gat), .ZN(new_n276_));
  INV_X1    g075(.A(G1gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT14), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT79), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(KEYINPUT79), .B(KEYINPUT14), .C1(new_n276_), .C2(new_n277_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G15gat), .B(G22gat), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT80), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT80), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n287_), .A3(new_n284_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G1gat), .B(G8gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n287_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n292_));
  AOI211_X1 g091(.A(KEYINPUT80), .B(new_n283_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n275_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G57gat), .B(G64gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT11), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G71gat), .B(G78gat), .Z(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(KEYINPUT11), .B2(new_n297_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n300_), .B(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n290_), .A2(new_n294_), .A3(new_n275_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n303_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n290_), .A2(new_n294_), .A3(new_n275_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(new_n295_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G127gat), .B(G155gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT16), .ZN(new_n310_));
  XOR2_X1   g109(.A(G183gat), .B(G211gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT17), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n305_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n308_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT17), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(KEYINPUT81), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT81), .B1(new_n315_), .B2(new_n317_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n314_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n315_), .A2(new_n317_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT81), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n318_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(KEYINPUT82), .A3(new_n314_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n274_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT13), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n332_), .A2(KEYINPUT71), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(KEYINPUT71), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n306_), .A2(KEYINPUT12), .A3(new_n245_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n254_), .A2(new_n303_), .A3(new_n255_), .ZN(new_n338_));
  INV_X1    g137(.A(G230gat), .ZN(new_n339_));
  INV_X1    g138(.A(G233gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n244_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n239_), .A2(new_n240_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n223_), .B2(KEYINPUT65), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n216_), .B1(new_n347_), .B2(new_n235_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n345_), .B1(new_n348_), .B2(new_n230_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT66), .B1(new_n349_), .B2(new_n229_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n255_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n306_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT12), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT69), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n303_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n355_), .A2(new_n356_), .A3(KEYINPUT12), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n337_), .B(new_n344_), .C1(new_n354_), .C2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n338_), .A2(KEYINPUT68), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n352_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n338_), .A2(KEYINPUT68), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n341_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G120gat), .B(G148gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT5), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G176gat), .B(G204gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n358_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n358_), .B2(new_n362_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT70), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n358_), .A2(new_n362_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n366_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT70), .B1(new_n374_), .B2(new_n368_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n334_), .B(new_n336_), .C1(new_n372_), .C2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n371_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(KEYINPUT70), .A3(new_n368_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT71), .A4(new_n332_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n376_), .A2(KEYINPUT72), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT72), .B1(new_n376_), .B2(new_n379_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n331_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(KEYINPUT83), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G141gat), .A2(G148gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(KEYINPUT91), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT2), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT91), .ZN(new_n390_));
  OAI22_X1  g189(.A1(new_n390_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n386_), .A2(new_n389_), .A3(new_n391_), .A4(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G155gat), .B(G162gat), .Z(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n384_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n396_), .A2(new_n387_), .ZN(new_n397_));
  INV_X1    g196(.A(G155gat), .ZN(new_n398_));
  INV_X1    g197(.A(G162gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT1), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT1), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(G155gat), .A3(G162gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n399_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n395_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT29), .ZN(new_n407_));
  NAND2_X1  g206(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(G233gat), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G211gat), .B(G218gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G197gat), .B(G204gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n412_), .B1(new_n414_), .B2(KEYINPUT21), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT21), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n413_), .B(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n417_), .B2(new_n412_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n407_), .A2(new_n411_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT94), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT94), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n407_), .A2(new_n418_), .A3(new_n421_), .A4(new_n411_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n411_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n393_), .A2(new_n394_), .B1(new_n397_), .B2(new_n404_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n418_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n420_), .A2(new_n422_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G78gat), .B(G106gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n420_), .A2(new_n422_), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n428_), .B(KEYINPUT96), .Z(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(new_n423_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G22gat), .B(G50gat), .Z(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n406_), .B2(KEYINPUT29), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n406_), .A2(KEYINPUT29), .A3(new_n435_), .ZN(new_n440_));
  OR3_X1    g239(.A1(new_n437_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n430_), .A2(KEYINPUT97), .A3(new_n434_), .A4(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT97), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n434_), .A2(new_n443_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n427_), .A2(new_n429_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n434_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n427_), .A2(new_n432_), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n443_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G183gat), .ZN(new_n456_));
  INV_X1    g255(.A(G190gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT23), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT23), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(G183gat), .A3(G190gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(KEYINPUT88), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n457_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n463_), .B(KEYINPUT23), .C1(new_n456_), .C2(new_n457_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(G169gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n469_));
  INV_X1    g268(.A(G169gat), .ZN(new_n470_));
  INV_X1    g269(.A(G176gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT87), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(G169gat), .B2(G176gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT24), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G169gat), .A2(G176gat), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n472_), .A2(new_n474_), .A3(KEYINPUT24), .A4(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT25), .B(G183gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT26), .B(G190gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n458_), .A2(new_n460_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n477_), .A2(new_n479_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n468_), .A2(new_n469_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n469_), .B1(new_n468_), .B2(new_n484_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n418_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n462_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n467_), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT98), .B(KEYINPUT24), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n475_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n491_), .A2(new_n464_), .A3(new_n482_), .A4(new_n461_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n472_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(new_n490_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n489_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n495_), .A2(new_n418_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n487_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G226gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT19), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n486_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n418_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n468_), .A2(new_n469_), .A3(new_n484_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT20), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n495_), .B2(new_n418_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n501_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G8gat), .B(G36gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT18), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT103), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n485_), .A2(new_n486_), .A3(new_n418_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n495_), .A2(new_n418_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT20), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n500_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n500_), .A2(new_n507_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n487_), .A2(new_n496_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n514_), .A3(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n516_), .A2(new_n517_), .A3(KEYINPUT27), .A4(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(KEYINPUT27), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n514_), .B1(new_n501_), .B2(new_n509_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT103), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n523_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n506_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n515_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n524_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT27), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n525_), .A2(new_n528_), .A3(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n455_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G127gat), .B(G134gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G113gat), .B(G120gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n538_), .A3(KEYINPUT90), .ZN(new_n542_));
  INV_X1    g341(.A(G127gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(G134gat), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n543_), .A2(G134gat), .ZN(new_n545_));
  INV_X1    g344(.A(G120gat), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n546_), .A2(G113gat), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(G113gat), .ZN(new_n548_));
  OAI22_X1  g347(.A1(new_n544_), .A2(new_n545_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n542_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(new_n424_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n539_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n552_), .A2(new_n395_), .A3(new_n405_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT4), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n406_), .A2(new_n541_), .A3(new_n542_), .A4(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT4), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G225gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n554_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n553_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n555_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n558_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G1gat), .B(G29gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT99), .B(G85gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT0), .B(G57gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n560_), .A2(new_n569_), .A3(new_n563_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n485_), .A2(new_n486_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G227gat), .A2(G233gat), .ZN(new_n576_));
  INV_X1    g375(.A(G15gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT30), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n575_), .B(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(new_n550_), .Z(new_n581_));
  XOR2_X1   g380(.A(G71gat), .B(G99gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(G43gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT31), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n580_), .B(new_n550_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n584_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n536_), .A2(new_n574_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n514_), .A2(KEYINPUT32), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n521_), .A2(new_n523_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT100), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT100), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n521_), .A2(new_n523_), .A3(new_n594_), .A4(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n591_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n510_), .A2(new_n597_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT102), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n569_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n559_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n569_), .B1(new_n562_), .B2(new_n558_), .ZN(new_n603_));
  OAI22_X1  g402(.A1(new_n601_), .A2(KEYINPUT33), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n601_), .A2(KEYINPUT33), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n532_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n596_), .A2(new_n598_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n448_), .A2(new_n444_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n525_), .A2(new_n528_), .A3(new_n534_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n573_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n610_), .A2(new_n611_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n590_), .B1(new_n614_), .B2(new_n589_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G169gat), .B(G197gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n290_), .A2(new_n294_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n256_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n621_), .A2(G229gat), .A3(G233gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT85), .Z(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n212_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT84), .B1(new_n620_), .B2(new_n256_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n212_), .A2(KEYINPUT84), .A3(new_n290_), .A4(new_n294_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n625_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n619_), .B1(new_n622_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n622_), .A2(new_n630_), .A3(new_n619_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT86), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n622_), .A2(new_n630_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n618_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT86), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n631_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n615_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n382_), .B2(KEYINPUT83), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n574_), .A2(G1gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n383_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n383_), .A2(new_n642_), .A3(KEYINPUT38), .A4(new_n643_), .ZN(new_n647_));
  AND4_X1   g446(.A1(new_n574_), .A2(new_n612_), .A3(new_n589_), .A4(new_n611_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n612_), .A2(new_n613_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n596_), .A2(new_n598_), .A3(new_n608_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n608_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n606_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n652_), .B2(new_n455_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n589_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n648_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n655_), .A2(new_n321_), .A3(new_n272_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n376_), .A2(KEYINPUT72), .A3(new_n379_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n376_), .A2(new_n379_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT72), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n632_), .A2(new_n633_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n656_), .A2(new_n657_), .A3(new_n660_), .A4(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n574_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n646_), .A2(new_n647_), .A3(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT104), .ZN(G1324gat));
  NAND2_X1  g465(.A1(new_n383_), .A2(new_n642_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n276_), .A3(new_n535_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n380_), .A2(new_n381_), .A3(new_n661_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n535_), .A3(new_n656_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n672_), .B2(G8gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n670_), .B(G8gat), .C1(new_n663_), .C2(new_n612_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(KEYINPUT106), .A2(KEYINPUT39), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .A4(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n675_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n677_), .B(new_n678_), .C1(new_n681_), .C2(new_n673_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n669_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n669_), .A2(new_n680_), .A3(KEYINPUT40), .A4(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  NAND3_X1  g486(.A1(new_n668_), .A2(new_n577_), .A3(new_n589_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n663_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n577_), .B1(new_n689_), .B2(new_n589_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n691_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n688_), .B1(new_n695_), .B2(new_n696_), .ZN(G1326gat));
  OAI21_X1  g496(.A(G22gat), .B1(new_n663_), .B2(new_n611_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT42), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n611_), .A2(G22gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n667_), .B2(new_n700_), .ZN(G1327gat));
  AOI21_X1  g500(.A(KEYINPUT82), .B1(new_n327_), .B2(new_n314_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n314_), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n322_), .B(new_n703_), .C1(new_n326_), .C2(new_n318_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n272_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n329_), .A2(KEYINPUT110), .A3(new_n272_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n653_), .A2(new_n654_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n639_), .B1(new_n710_), .B2(new_n590_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n709_), .A2(new_n660_), .A3(new_n711_), .A4(new_n657_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n713_), .B2(new_n573_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n329_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n270_), .A2(KEYINPUT37), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n272_), .A2(new_n273_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n655_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n615_), .A2(new_n720_), .A3(new_n274_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n715_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n671_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT44), .B1(new_n723_), .B2(KEYINPUT109), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n725_), .B(new_n726_), .C1(new_n722_), .C2(new_n671_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n573_), .A2(G29gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n714_), .B1(new_n729_), .B2(new_n730_), .ZN(G1328gat));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT111), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n612_), .A2(G36gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n713_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n735_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n712_), .A2(KEYINPUT45), .A3(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n733_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n535_), .B1(new_n724_), .B2(new_n727_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(G36gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n732_), .A2(KEYINPUT111), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n742_), .B(new_n739_), .C1(new_n740_), .C2(G36gat), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1329gat));
  NAND2_X1  g545(.A1(new_n589_), .A2(G43gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n712_), .A2(new_n654_), .ZN(new_n748_));
  OAI22_X1  g547(.A1(new_n728_), .A2(new_n747_), .B1(G43gat), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g549(.A(G50gat), .B1(new_n713_), .B2(new_n455_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n455_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n729_), .B2(new_n752_), .ZN(G1331gat));
  AOI21_X1  g552(.A(new_n662_), .B1(new_n660_), .B2(new_n657_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n615_), .ZN(new_n755_));
  OR4_X1    g554(.A1(G57gat), .A2(new_n755_), .A3(new_n331_), .A4(new_n574_), .ZN(new_n756_));
  NOR4_X1   g555(.A1(new_n655_), .A2(new_n640_), .A3(new_n329_), .A4(new_n272_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n380_), .A2(new_n381_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G57gat), .B1(new_n760_), .B2(new_n574_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(new_n761_), .ZN(G1332gat));
  OR4_X1    g561(.A1(G64gat), .A2(new_n755_), .A3(new_n331_), .A4(new_n612_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n535_), .A3(new_n757_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(G64gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n764_), .B2(G64gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1333gat));
  OR4_X1    g567(.A1(G71gat), .A2(new_n755_), .A3(new_n331_), .A4(new_n654_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n759_), .A2(new_n589_), .A3(new_n757_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(G71gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G71gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1334gat));
  OR4_X1    g573(.A1(G78gat), .A2(new_n755_), .A3(new_n331_), .A4(new_n611_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n759_), .A2(new_n455_), .A3(new_n757_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G78gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G78gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1335gat));
  INV_X1    g579(.A(new_n754_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(new_n715_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n655_), .A2(new_n718_), .A3(KEYINPUT43), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n720_), .B1(new_n615_), .B2(new_n274_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(KEYINPUT112), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G85gat), .B1(new_n788_), .B2(new_n574_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT110), .B1(new_n329_), .B2(new_n272_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n706_), .B(new_n271_), .C1(new_n323_), .C2(new_n328_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n755_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n213_), .A3(new_n573_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n789_), .A2(new_n794_), .ZN(G1336gat));
  AOI21_X1  g594(.A(G92gat), .B1(new_n793_), .B2(new_n535_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n788_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n535_), .A2(G92gat), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT113), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n797_), .B2(new_n799_), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n788_), .B2(new_n654_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n654_), .A2(new_n228_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n793_), .A2(new_n802_), .B1(new_n803_), .B2(KEYINPUT51), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n803_), .A2(KEYINPUT51), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n805_), .B(new_n807_), .ZN(G1338gat));
  NAND3_X1  g607(.A1(new_n793_), .A2(new_n238_), .A3(new_n455_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n722_), .A2(KEYINPUT115), .A3(new_n455_), .A4(new_n754_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n811_), .A2(G106gat), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n329_), .B(new_n455_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n781_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n810_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  AND4_X1   g615(.A1(new_n810_), .A2(new_n815_), .A3(G106gat), .A4(new_n811_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n809_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT53), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n809_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1339gat));
  NAND3_X1  g621(.A1(new_n536_), .A2(new_n573_), .A3(new_n589_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n337_), .B(new_n338_), .C1(new_n354_), .C2(new_n357_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n341_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n337_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n352_), .A2(KEYINPUT69), .A3(new_n353_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n356_), .B1(new_n355_), .B2(KEYINPUT12), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT117), .B1(new_n830_), .B2(new_n344_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n826_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n358_), .A2(new_n834_), .A3(new_n832_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT56), .B(new_n366_), .C1(new_n833_), .C2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n358_), .A2(new_n834_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n839_), .A2(KEYINPUT55), .B1(new_n341_), .B2(new_n825_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n367_), .B1(new_n840_), .B2(new_n835_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT119), .B1(new_n841_), .B2(KEYINPUT56), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n366_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n838_), .B1(new_n842_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n628_), .A2(new_n629_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n625_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n618_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n633_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n368_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n824_), .B1(new_n847_), .B2(new_n852_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n827_), .B(new_n343_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT55), .B1(new_n854_), .B2(KEYINPUT117), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n835_), .A3(new_n826_), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT119), .B(KEYINPUT56), .C1(new_n856_), .C2(new_n366_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n844_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n837_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n852_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(KEYINPUT58), .A3(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n853_), .A2(new_n861_), .A3(new_n274_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n856_), .A2(new_n864_), .A3(KEYINPUT56), .A4(new_n366_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n369_), .B1(new_n636_), .B2(new_n631_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n837_), .A2(KEYINPUT118), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT56), .B1(new_n856_), .B2(new_n366_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n865_), .B(new_n866_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n851_), .A2(new_n378_), .A3(new_n377_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n863_), .B1(new_n872_), .B2(new_n271_), .ZN(new_n873_));
  AOI211_X1 g672(.A(KEYINPUT57), .B(new_n272_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n862_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n321_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n718_), .A2(new_n715_), .A3(new_n639_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n878_));
  OR3_X1    g677(.A1(new_n877_), .A2(new_n658_), .A3(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n877_), .B2(new_n658_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n823_), .B1(new_n876_), .B2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(G113gat), .B1(new_n883_), .B2(new_n662_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n843_), .A2(new_n845_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(KEYINPUT118), .A3(new_n837_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n865_), .A2(new_n866_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n870_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT57), .B1(new_n888_), .B2(new_n272_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n872_), .A2(new_n863_), .A3(new_n271_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n715_), .B1(new_n891_), .B2(new_n862_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(new_n881_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n823_), .A2(KEYINPUT59), .ZN(new_n894_));
  INV_X1    g693(.A(new_n823_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n321_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n891_), .B2(new_n862_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n897_), .B2(new_n881_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n893_), .A2(new_n894_), .B1(new_n898_), .B2(KEYINPUT59), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT120), .B(G113gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n640_), .A2(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT121), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n884_), .B1(new_n899_), .B2(new_n902_), .ZN(G1340gat));
  OAI21_X1  g702(.A(new_n894_), .B1(new_n892_), .B2(new_n881_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n759_), .B(new_n904_), .C1(new_n883_), .C2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(G120gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n546_), .B1(new_n758_), .B2(KEYINPUT60), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n883_), .B(new_n908_), .C1(KEYINPUT60), .C2(new_n546_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1341gat));
  OAI211_X1 g709(.A(new_n715_), .B(new_n895_), .C1(new_n897_), .C2(new_n881_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n543_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT122), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n321_), .A2(new_n543_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n904_), .B(new_n914_), .C1(new_n883_), .C2(new_n905_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n911_), .A2(new_n916_), .A3(new_n543_), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n913_), .A2(new_n915_), .A3(new_n917_), .ZN(G1342gat));
  AOI21_X1  g717(.A(G134gat), .B1(new_n883_), .B2(new_n272_), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT123), .B(G134gat), .Z(new_n920_));
  NOR2_X1   g719(.A1(new_n718_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n899_), .B2(new_n921_), .ZN(G1343gat));
  NAND2_X1  g721(.A1(new_n876_), .A2(new_n882_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n589_), .A2(new_n535_), .A3(new_n611_), .A4(new_n574_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n923_), .A2(new_n662_), .A3(new_n924_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT124), .B(G141gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1344gat));
  NAND3_X1  g726(.A1(new_n923_), .A2(new_n759_), .A3(new_n924_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g728(.A1(new_n923_), .A2(new_n715_), .A3(new_n924_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT61), .B(G155gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n930_), .B(new_n931_), .ZN(G1346gat));
  NAND2_X1  g731(.A1(new_n923_), .A2(new_n924_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G162gat), .B1(new_n933_), .B2(new_n718_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n272_), .A2(new_n399_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n933_), .B2(new_n935_), .ZN(G1347gat));
  NOR4_X1   g735(.A1(new_n654_), .A2(new_n612_), .A3(new_n573_), .A4(new_n455_), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n662_), .B(new_n937_), .C1(new_n892_), .C2(new_n881_), .ZN(new_n938_));
  OAI21_X1  g737(.A(KEYINPUT62), .B1(new_n938_), .B2(KEYINPUT22), .ZN(new_n939_));
  OAI21_X1  g738(.A(G169gat), .B1(new_n938_), .B2(KEYINPUT62), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  OAI211_X1 g740(.A(KEYINPUT62), .B(G169gat), .C1(new_n938_), .C2(KEYINPUT22), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1348gat));
  NAND3_X1  g742(.A1(new_n893_), .A2(new_n759_), .A3(new_n937_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n923_), .A2(new_n937_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n758_), .A2(new_n471_), .ZN(new_n946_));
  AOI22_X1  g745(.A1(new_n471_), .A2(new_n944_), .B1(new_n945_), .B2(new_n946_), .ZN(G1349gat));
  NAND2_X1  g746(.A1(new_n893_), .A2(new_n937_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n321_), .A2(new_n480_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n923_), .A2(new_n715_), .A3(new_n937_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n949_), .A2(new_n950_), .B1(new_n951_), .B2(new_n456_), .ZN(G1350gat));
  OAI211_X1 g751(.A(new_n274_), .B(new_n937_), .C1(new_n892_), .C2(new_n881_), .ZN(new_n953_));
  AND3_X1   g752(.A1(new_n953_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n954_));
  AOI21_X1  g753(.A(KEYINPUT125), .B1(new_n953_), .B2(G190gat), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n272_), .A2(new_n481_), .ZN(new_n956_));
  OAI22_X1  g755(.A1(new_n954_), .A2(new_n955_), .B1(new_n948_), .B2(new_n956_), .ZN(G1351gat));
  NAND3_X1  g756(.A1(new_n654_), .A2(new_n613_), .A3(new_n535_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n958_), .B1(new_n876_), .B2(new_n882_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(new_n662_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(KEYINPUT126), .B(G197gat), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n960_), .B(new_n961_), .ZN(G1352gat));
  NAND2_X1  g761(.A1(new_n959_), .A2(new_n759_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g763(.A(new_n321_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n959_), .A2(new_n965_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  OR2_X1    g766(.A1(new_n967_), .A2(KEYINPUT127), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(KEYINPUT127), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n966_), .A2(new_n968_), .A3(new_n969_), .ZN(new_n970_));
  NAND4_X1  g769(.A1(new_n959_), .A2(KEYINPUT127), .A3(new_n965_), .A4(new_n967_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(G1354gat));
  INV_X1    g771(.A(G218gat), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n959_), .A2(new_n973_), .A3(new_n272_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n959_), .A2(new_n274_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n975_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n974_), .B1(new_n976_), .B2(new_n973_), .ZN(G1355gat));
endmodule


