//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(G113gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G120gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G227gat), .A2(G233gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT30), .Z(new_n210_));
  XNOR2_X1  g009(.A(new_n208_), .B(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G71gat), .B(G99gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT31), .ZN(new_n213_));
  XOR2_X1   g012(.A(G15gat), .B(G43gat), .Z(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(G183gat), .B2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT22), .B(G169gat), .Z(new_n223_));
  OAI211_X1 g022(.A(new_n221_), .B(new_n222_), .C1(G176gat), .C2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT81), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n219_), .A3(new_n218_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT81), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n226_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G183gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT25), .B(G183gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n235_), .B(new_n239_), .C1(new_n240_), .C2(new_n238_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n229_), .A2(new_n231_), .A3(new_n234_), .A4(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n224_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n215_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n211_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n211_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT18), .B(G64gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G92gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G8gat), .B(G36gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT94), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT91), .Z(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT19), .Z(new_n258_));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n240_), .A2(KEYINPUT92), .ZN(new_n260_));
  INV_X1    g059(.A(G183gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT25), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n237_), .A2(new_n262_), .A3(KEYINPUT92), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n235_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n232_), .A2(KEYINPUT93), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n232_), .A2(KEYINPUT93), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n233_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n230_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n224_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT21), .ZN(new_n271_));
  INV_X1    g070(.A(G197gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(G204gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT88), .ZN(new_n274_));
  INV_X1    g073(.A(G204gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n274_), .B1(new_n275_), .B2(G197gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT89), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n271_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G211gat), .B(G218gat), .Z(new_n281_));
  OAI211_X1 g080(.A(new_n280_), .B(new_n281_), .C1(new_n279_), .C2(new_n278_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n278_), .B2(new_n271_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n275_), .A2(G197gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n272_), .A2(G204gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n271_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n286_), .A2(KEYINPUT87), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(KEYINPUT87), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n259_), .B1(new_n270_), .B2(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n282_), .A2(new_n224_), .A3(new_n289_), .A4(new_n242_), .ZN(new_n292_));
  AOI211_X1 g091(.A(new_n255_), .B(new_n258_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n270_), .A2(new_n290_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(KEYINPUT20), .A3(new_n292_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n258_), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT94), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n290_), .A2(new_n243_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n269_), .A2(new_n282_), .A3(new_n289_), .A4(new_n224_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(KEYINPUT20), .A3(new_n300_), .A4(new_n258_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT95), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n254_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n295_), .A2(new_n296_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n255_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n295_), .A2(KEYINPUT94), .A3(new_n296_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT95), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n301_), .B(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n253_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT96), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n303_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n307_), .A2(new_n309_), .A3(KEYINPUT96), .A4(new_n253_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT0), .B(G57gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(G85gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(G1gat), .B(G29gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G155gat), .ZN(new_n319_));
  INV_X1    g118(.A(G162gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n319_), .A2(new_n320_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT85), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n323_), .ZN(new_n327_));
  OAI211_X1 g126(.A(KEYINPUT85), .B(new_n321_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT84), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n322_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335_));
  INV_X1    g134(.A(G141gat), .ZN(new_n336_));
  INV_X1    g135(.A(G148gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n330_), .A2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .A4(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n343_), .A2(KEYINPUT86), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(KEYINPUT86), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n334_), .B(new_n321_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n333_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n204_), .B(G120gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n206_), .A2(new_n333_), .A3(new_n346_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n318_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT98), .Z(new_n355_));
  NAND3_X1  g154(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT4), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(KEYINPUT4), .B2(new_n349_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n355_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(new_n353_), .C1(KEYINPUT4), .C2(new_n349_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n351_), .A2(new_n352_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n318_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT33), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n361_), .A2(KEYINPUT97), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n361_), .B2(KEYINPUT97), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n314_), .A2(new_n358_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n359_), .A2(new_n360_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n318_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n361_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n253_), .A2(KEYINPUT32), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n295_), .A2(new_n296_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n259_), .B1(new_n290_), .B2(new_n243_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n258_), .B1(new_n373_), .B2(new_n300_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n371_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n307_), .A2(new_n309_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n370_), .B(new_n375_), .C1(new_n371_), .C2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n249_), .B1(new_n366_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT90), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n347_), .A2(KEYINPUT29), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n290_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n333_), .B2(new_n346_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n290_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G78gat), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n382_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n388_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n390_));
  INV_X1    g189(.A(G106gat), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n381_), .B1(new_n380_), .B2(new_n290_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n385_), .A2(new_n386_), .A3(new_n383_), .ZN(new_n394_));
  OAI21_X1  g193(.A(G78gat), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n382_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n396_));
  AOI21_X1  g195(.A(G106gat), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n379_), .B1(new_n392_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n333_), .A2(new_n346_), .A3(new_n384_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G22gat), .B(G50gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT28), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n399_), .B(new_n401_), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n391_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n395_), .A2(G106gat), .A3(new_n396_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(KEYINPUT90), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n398_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n379_), .B(new_n402_), .C1(new_n392_), .C2(new_n397_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n378_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT27), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n312_), .A2(new_n411_), .A3(new_n313_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n254_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n310_), .A2(KEYINPUT27), .A3(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n370_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n369_), .A2(KEYINPUT99), .A3(new_n361_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n407_), .A2(new_n408_), .A3(new_n248_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n248_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n415_), .B(new_n420_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n410_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G43gat), .B(G50gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G29gat), .B(G36gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n427_), .B(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G15gat), .B(G22gat), .ZN(new_n431_));
  INV_X1    g230(.A(G1gat), .ZN(new_n432_));
  INV_X1    g231(.A(G8gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT14), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G1gat), .B(G8gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n430_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n427_), .B(new_n428_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT15), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n430_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n438_), .B1(new_n443_), .B2(new_n437_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G229gat), .A2(G233gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n439_), .B(new_n437_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G113gat), .B(G141gat), .ZN(new_n449_));
  INV_X1    g248(.A(G169gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(new_n272_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n448_), .B(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G85gat), .A2(G92gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(KEYINPUT9), .ZN(new_n457_));
  INV_X1    g256(.A(G99gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT10), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT10), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(G99gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n391_), .A2(KEYINPUT64), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT64), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n457_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n468_));
  AND3_X1   g267(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G99gat), .A2(G106gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(KEYINPUT65), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G85gat), .ZN(new_n478_));
  INV_X1    g277(.A(G92gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(KEYINPUT9), .A3(new_n456_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n467_), .A2(new_n477_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(G57gat), .ZN(new_n484_));
  INV_X1    g283(.A(G64gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G57gat), .A2(G64gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G71gat), .B(G78gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT11), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n486_), .A2(new_n492_), .A3(new_n487_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n488_), .A2(new_n490_), .A3(KEYINPUT11), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n458_), .A2(new_n391_), .A3(KEYINPUT67), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT66), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n498_), .A3(KEYINPUT7), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n469_), .A2(new_n470_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501_));
  NOR2_X1   g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(KEYINPUT66), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT66), .B1(new_n502_), .B2(KEYINPUT67), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n499_), .B(new_n500_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n480_), .A2(new_n456_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT68), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n480_), .A2(new_n508_), .A3(new_n456_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT8), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT8), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n471_), .A2(new_n476_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n499_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n513_), .B(new_n510_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n516_));
  AOI211_X1 g315(.A(new_n483_), .B(new_n496_), .C1(new_n512_), .C2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n513_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n515_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT8), .B1(new_n519_), .B2(new_n477_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n520_), .B2(new_n510_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n496_), .B1(new_n521_), .B2(new_n483_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n517_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n496_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(new_n523_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n512_), .A2(new_n516_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n482_), .A2(KEYINPUT70), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n467_), .A2(new_n477_), .A3(new_n529_), .A4(new_n481_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n527_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n527_), .B2(new_n531_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n526_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G230gat), .A2(G233gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n524_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n525_), .B1(new_n527_), .B2(new_n482_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n517_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n455_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n540_), .A2(new_n455_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G120gat), .B(G148gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n275_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT5), .ZN(new_n545_));
  INV_X1    g344(.A(G176gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OR3_X1    g347(.A1(new_n541_), .A2(new_n542_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n548_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT13), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT72), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n549_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(KEYINPUT72), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n549_), .A2(new_n550_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT73), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n549_), .A2(new_n550_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n554_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n549_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n454_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n443_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n521_), .A2(new_n483_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n439_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT34), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT35), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n568_), .A2(KEYINPUT35), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n564_), .A2(new_n566_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT76), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n527_), .A2(new_n531_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT71), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n527_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n578_), .A2(new_n443_), .B1(new_n439_), .B2(new_n565_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n573_), .B(new_n574_), .C1(new_n579_), .C2(new_n569_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(KEYINPUT76), .A3(new_n572_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(G134gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n320_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(KEYINPUT36), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT78), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT77), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n585_), .B(KEYINPUT36), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n580_), .A2(new_n590_), .A3(new_n591_), .A4(new_n581_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT77), .B1(new_n589_), .B2(KEYINPUT37), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n580_), .A2(new_n581_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n597_), .B2(new_n591_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n588_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n437_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n496_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT79), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT16), .B(G183gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G211gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n603_), .B(new_n609_), .Z(new_n610_));
  INV_X1    g409(.A(new_n602_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n608_), .A3(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n595_), .A2(new_n599_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n424_), .A2(new_n563_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n432_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n420_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT100), .Z(new_n620_));
  OAI21_X1  g419(.A(new_n618_), .B1(new_n617_), .B2(new_n420_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT101), .Z(new_n622_));
  NAND2_X1  g421(.A1(new_n409_), .A2(new_n249_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n407_), .A2(new_n408_), .A3(new_n248_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n419_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n625_), .A2(new_n415_), .B1(new_n378_), .B2(new_n409_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n588_), .A2(new_n592_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n597_), .A2(new_n591_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT77), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n613_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n626_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n563_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n634_), .B2(new_n420_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n620_), .A2(new_n622_), .A3(new_n635_), .ZN(G1324gat));
  INV_X1    g435(.A(new_n415_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n616_), .A2(new_n433_), .A3(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G8gat), .B1(new_n634_), .B2(new_n415_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(KEYINPUT39), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(KEYINPUT39), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n616_), .A2(new_n645_), .A3(new_n249_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G15gat), .B1(new_n634_), .B2(new_n248_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n409_), .B(KEYINPUT102), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n616_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G22gat), .B1(new_n634_), .B2(new_n655_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT103), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT103), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n657_), .A2(KEYINPUT42), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT42), .B1(new_n657_), .B2(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n654_), .B1(new_n659_), .B2(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n593_), .A2(new_n594_), .B1(new_n598_), .B2(new_n588_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n424_), .B2(new_n664_), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT43), .B(new_n663_), .C1(new_n410_), .C2(new_n423_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n563_), .B(new_n632_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT43), .B1(new_n626_), .B2(new_n663_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n424_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n563_), .A4(new_n632_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n673_), .A3(new_n419_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G29gat), .ZN(new_n675_));
  AND4_X1   g474(.A1(new_n563_), .A2(new_n424_), .A3(new_n631_), .A4(new_n632_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n420_), .A2(G29gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT104), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n677_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(KEYINPUT105), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(KEYINPUT105), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n669_), .A2(new_n673_), .A3(new_n637_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n676_), .A2(new_n686_), .A3(new_n637_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT45), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n682_), .B(new_n683_), .C1(new_n685_), .C2(new_n688_), .ZN(new_n689_));
  AND4_X1   g488(.A1(KEYINPUT105), .A2(new_n685_), .A3(new_n681_), .A4(new_n688_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1329gat));
  INV_X1    g490(.A(G43gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n248_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n669_), .A2(new_n673_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n692_), .B1(new_n677_), .B2(new_n248_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n695_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n694_), .A2(new_n696_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT106), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT47), .B1(new_n703_), .B2(new_n697_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1330gat));
  INV_X1    g504(.A(new_n409_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n669_), .A2(new_n673_), .A3(new_n706_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n707_), .A2(KEYINPUT107), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(KEYINPUT107), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(G50gat), .A3(new_n709_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n655_), .A2(G50gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n677_), .B2(new_n711_), .ZN(G1331gat));
  NAND2_X1  g511(.A1(new_n556_), .A2(new_n562_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n453_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n424_), .A3(new_n615_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n419_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n633_), .A2(new_n714_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(new_n420_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n719_), .B2(G57gat), .ZN(G1332gat));
  NAND3_X1  g519(.A1(new_n716_), .A2(new_n485_), .A3(new_n637_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G64gat), .B1(new_n718_), .B2(new_n415_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT48), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(KEYINPUT48), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(G1333gat));
  OAI21_X1  g524(.A(G71gat), .B1(new_n718_), .B2(new_n248_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT49), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(KEYINPUT49), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n248_), .A2(G71gat), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT108), .Z(new_n730_));
  OAI22_X1  g529(.A1(new_n727_), .A2(new_n728_), .B1(new_n715_), .B2(new_n730_), .ZN(G1334gat));
  NAND3_X1  g530(.A1(new_n633_), .A2(new_n653_), .A3(new_n714_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G78gat), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT109), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(KEYINPUT109), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736_));
  OR3_X1    g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n716_), .A2(new_n388_), .A3(new_n653_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(G1335gat));
  NOR3_X1   g539(.A1(new_n713_), .A2(new_n453_), .A3(new_n613_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n741_), .A2(new_n424_), .A3(new_n631_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n478_), .A3(new_n419_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n672_), .A2(new_n741_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(new_n419_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n745_), .B2(new_n478_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT110), .Z(G1336gat));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n637_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n742_), .A2(new_n479_), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n748_), .A2(G92gat), .B1(new_n637_), .B2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT111), .Z(G1337gat));
  NAND3_X1  g550(.A1(new_n742_), .A2(new_n462_), .A3(new_n249_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT112), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n458_), .B1(new_n744_), .B2(new_n249_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n742_), .A2(new_n466_), .A3(new_n706_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n672_), .A2(new_n706_), .A3(new_n741_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(G106gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G106gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g563(.A1(new_n637_), .A2(new_n420_), .A3(new_n623_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n526_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n527_), .A2(new_n482_), .A3(new_n525_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n539_), .B2(KEYINPUT12), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n767_), .A2(new_n769_), .A3(new_n538_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n538_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(KEYINPUT55), .B2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n524_), .A2(new_n535_), .A3(KEYINPUT55), .A4(new_n536_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n548_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT114), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n536_), .B1(new_n524_), .B2(new_n535_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n537_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n547_), .B1(new_n780_), .B2(new_n773_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT56), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n781_), .B2(KEYINPUT56), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n777_), .A2(new_n782_), .A3(new_n784_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n448_), .A2(new_n452_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n445_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n444_), .A2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n788_), .B(new_n452_), .C1(new_n787_), .C2(new_n447_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n549_), .A2(new_n786_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n785_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n664_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n785_), .A2(KEYINPUT58), .A3(new_n790_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT58), .B1(new_n785_), .B2(new_n790_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT115), .B1(new_n797_), .B2(new_n663_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n781_), .A2(KEYINPUT56), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n781_), .A2(KEYINPUT56), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n453_), .B(new_n549_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n557_), .A2(new_n786_), .A3(new_n789_), .ZN(new_n804_));
  AOI221_X4 g603(.A(new_n800_), .B1(new_n627_), .B2(new_n629_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n804_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT57), .B1(new_n806_), .B2(new_n630_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n613_), .B1(new_n799_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n454_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT113), .B1(new_n614_), .B2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n453_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n663_), .A4(new_n613_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n811_), .A2(new_n814_), .A3(KEYINPUT54), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT54), .B1(new_n811_), .B2(new_n814_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n765_), .B1(new_n809_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(G113gat), .B1(new_n819_), .B2(new_n453_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822_));
  OAI22_X1  g621(.A1(new_n809_), .A2(new_n822_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n823_));
  AOI211_X1 g622(.A(KEYINPUT117), .B(new_n613_), .C1(new_n799_), .C2(new_n808_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n821_), .B(new_n765_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n818_), .A2(new_n826_), .A3(KEYINPUT59), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n818_), .B2(KEYINPUT59), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n453_), .B(new_n825_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n820_), .B1(new_n830_), .B2(G113gat), .ZN(G1340gat));
  XNOR2_X1  g630(.A(KEYINPUT118), .B(G120gat), .ZN(new_n832_));
  INV_X1    g631(.A(new_n713_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n832_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT60), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n818_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT60), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n832_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n825_), .B(new_n836_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n841_), .B2(new_n833_), .ZN(G1341gat));
  AOI21_X1  g641(.A(G127gat), .B1(new_n819_), .B2(new_n613_), .ZN(new_n843_));
  OR2_X1    g642(.A1(KEYINPUT119), .A2(G127gat), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n825_), .B(new_n844_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(G127gat), .B1(new_n632_), .B2(KEYINPUT119), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n843_), .B1(new_n846_), .B2(new_n847_), .ZN(G1342gat));
  INV_X1    g647(.A(G134gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n663_), .A2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n825_), .B(new_n850_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n849_), .B1(new_n818_), .B2(new_n630_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT120), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1343gat));
  NOR2_X1   g654(.A1(new_n809_), .A2(new_n817_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n624_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n637_), .A2(new_n420_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n454_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT121), .B(G141gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1344gat));
  NOR2_X1   g661(.A1(new_n859_), .A2(new_n713_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(new_n337_), .ZN(G1345gat));
  NOR2_X1   g663(.A1(new_n859_), .A2(new_n632_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT61), .B(G155gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  NOR3_X1   g666(.A1(new_n859_), .A2(new_n320_), .A3(new_n663_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n857_), .A2(new_n631_), .A3(new_n858_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n320_), .B2(new_n869_), .ZN(G1347gat));
  NOR3_X1   g669(.A1(new_n415_), .A2(new_n419_), .A3(new_n248_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(KEYINPUT122), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n415_), .A2(new_n419_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(KEYINPUT122), .A3(new_n249_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n653_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n453_), .B(new_n875_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(G169gat), .A3(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n879_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n876_), .A2(G169gat), .A3(new_n881_), .A4(new_n877_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n880_), .B(new_n882_), .C1(new_n223_), .C2(new_n876_), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n856_), .A2(new_n706_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n872_), .A2(new_n874_), .ZN(new_n885_));
  AND4_X1   g684(.A1(G176gat), .A2(new_n884_), .A3(new_n833_), .A4(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n833_), .B(new_n875_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n889_), .B2(G176gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(KEYINPUT124), .A3(new_n546_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n886_), .B1(new_n890_), .B2(new_n891_), .ZN(G1349gat));
  OR2_X1    g691(.A1(new_n823_), .A2(new_n824_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n893_), .A2(new_n875_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n632_), .A2(new_n260_), .A3(new_n263_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n884_), .A2(new_n613_), .A3(new_n885_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n894_), .A2(new_n895_), .B1(new_n261_), .B2(new_n896_), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n235_), .A3(new_n631_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n893_), .A2(new_n664_), .A3(new_n875_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G190gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1351gat));
  OAI211_X1 g700(.A(new_n421_), .B(new_n873_), .C1(new_n809_), .C2(new_n817_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n454_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n272_), .ZN(G1352gat));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n713_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n905_), .B2(new_n906_), .ZN(G1353gat));
  NOR2_X1   g708(.A1(new_n902_), .A2(new_n632_), .ZN(new_n910_));
  OR2_X1    g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n910_), .A2(KEYINPUT126), .A3(new_n911_), .A4(new_n912_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  OR3_X1    g716(.A1(new_n910_), .A2(new_n917_), .A3(new_n911_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n915_), .A2(new_n916_), .B1(new_n918_), .B2(new_n919_), .ZN(G1354gat));
  INV_X1    g719(.A(G218gat), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n902_), .A2(new_n921_), .A3(new_n663_), .ZN(new_n922_));
  OR2_X1    g721(.A1(new_n902_), .A2(new_n630_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n921_), .B2(new_n923_), .ZN(G1355gat));
endmodule


