//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT82), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT82), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G155gat), .A3(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT83), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n206_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT1), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT83), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n204_), .A2(new_n206_), .A3(new_n212_), .A4(new_n207_), .ZN(new_n213_));
  OR2_X1    g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n209_), .A2(new_n211_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G141gat), .B(G148gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n205_), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n203_), .A2(KEYINPUT82), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n214_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n210_), .A2(KEYINPUT86), .A3(new_n214_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT85), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n229_), .A2(KEYINPUT84), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT84), .B1(new_n229_), .B2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n228_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n222_), .B(new_n223_), .C1(new_n225_), .C2(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n217_), .A2(new_n234_), .A3(KEYINPUT87), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT87), .B1(new_n217_), .B2(new_n234_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n202_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT28), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT28), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n239_), .B(new_n202_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G22gat), .B(G50gat), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n238_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G197gat), .B(G204gat), .Z(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT21), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G197gat), .B(G204gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT21), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G211gat), .B(G218gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  OR3_X1    g050(.A1(new_n247_), .A2(new_n250_), .A3(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n217_), .A2(new_n234_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n256_));
  OAI21_X1  g055(.A(new_n253_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(G228gat), .A3(G233gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n217_), .A2(new_n234_), .A3(KEYINPUT87), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT29), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G228gat), .A2(G233gat), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n253_), .A2(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n262_), .A2(KEYINPUT88), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT88), .B1(new_n262_), .B2(new_n264_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n258_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G78gat), .B(G106gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n258_), .B(new_n270_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n244_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT90), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT88), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n235_), .A2(new_n236_), .A3(new_n202_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n264_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n262_), .A2(KEYINPUT88), .A3(new_n264_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n280_), .A2(KEYINPUT90), .A3(new_n258_), .A4(new_n270_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n274_), .A2(new_n269_), .A3(new_n281_), .A4(new_n244_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT91), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n270_), .B1(new_n280_), .B2(new_n258_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n238_), .A2(new_n240_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n241_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n238_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT91), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n281_), .A4(new_n274_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n272_), .B1(new_n283_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT23), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(G176gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT24), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(KEYINPUT24), .A3(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n295_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n303_));
  INV_X1    g102(.A(G183gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT76), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G183gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n303_), .B1(new_n308_), .B2(KEYINPUT25), .ZN(new_n309_));
  INV_X1    g108(.A(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT26), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT26), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT77), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT77), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n316_), .B(new_n317_), .C1(new_n319_), .C2(new_n303_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n302_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n294_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT76), .B(G183gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n310_), .B2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(new_n296_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT78), .B1(new_n321_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n302_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n320_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n303_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(new_n324_), .B2(new_n318_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n316_), .B1(new_n333_), .B2(new_n317_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n330_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n325_), .A2(new_n327_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n253_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n329_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT20), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT94), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n344_), .B(new_n295_), .C1(new_n298_), .C2(new_n343_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n311_), .A2(new_n313_), .A3(KEYINPUT92), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT92), .B1(new_n311_), .B2(new_n313_), .ZN(new_n347_));
  XOR2_X1   g146(.A(KEYINPUT25), .B(G183gat), .Z(new_n348_));
  NOR3_X1   g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n342_), .B1(new_n345_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n347_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n317_), .A2(KEYINPUT92), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n343_), .A2(new_n298_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(new_n323_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n354_), .A2(new_n356_), .A3(KEYINPUT94), .A4(new_n344_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n295_), .B1(G183gat), .B2(G190gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n300_), .B(KEYINPUT95), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT22), .B(G169gat), .Z(new_n360_));
  OAI211_X1 g159(.A(new_n358_), .B(new_n359_), .C1(G176gat), .C2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n350_), .A2(new_n357_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n341_), .B1(new_n362_), .B2(new_n253_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n340_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT19), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n329_), .A2(new_n338_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n253_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n339_), .A2(new_n350_), .A3(new_n357_), .A4(new_n361_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n366_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n370_), .A2(KEYINPUT20), .A3(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n372_), .A3(KEYINPUT96), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT18), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  INV_X1    g177(.A(KEYINPUT96), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n339_), .B1(new_n329_), .B2(new_n338_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n370_), .A2(KEYINPUT20), .A3(new_n371_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n374_), .A2(KEYINPUT99), .A3(new_n378_), .A4(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n339_), .A2(new_n361_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n345_), .A2(new_n349_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT20), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n366_), .B1(new_n380_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT98), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT98), .B(new_n366_), .C1(new_n380_), .C2(new_n386_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n340_), .A2(new_n371_), .A3(new_n363_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n378_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n367_), .A2(new_n373_), .A3(new_n378_), .A4(new_n382_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT99), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n383_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT27), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n367_), .A2(new_n373_), .A3(new_n382_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n393_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n395_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(KEYINPUT27), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n399_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  INV_X1    g205(.A(G15gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT30), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G71gat), .B(G99gat), .ZN(new_n411_));
  INV_X1    g210(.A(G43gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n368_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n368_), .A2(new_n413_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n410_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n368_), .A2(new_n413_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n409_), .A3(new_n414_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT81), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G127gat), .B(G134gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G120gat), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n424_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n424_), .A3(KEYINPUT79), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT80), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT31), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n417_), .A2(new_n419_), .A3(KEYINPUT81), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n422_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n420_), .A2(new_n421_), .A3(new_n432_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n260_), .A2(new_n261_), .A3(new_n430_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n425_), .A2(new_n427_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n255_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(KEYINPUT4), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT97), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT97), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n438_), .A2(new_n443_), .A3(KEYINPUT4), .A4(new_n440_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n260_), .A2(new_n446_), .A3(new_n261_), .A4(new_n430_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G225gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n438_), .A2(new_n440_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(new_n449_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G29gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(G85gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT0), .B(G57gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n457_), .B(new_n458_), .Z(new_n459_));
  NAND3_X1  g258(.A1(new_n452_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n450_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n461_), .B1(new_n462_), .B2(new_n454_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n437_), .A2(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n293_), .A2(new_n405_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n437_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n283_), .A2(new_n292_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n272_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n464_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n392_), .A2(new_n393_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n473_), .B2(new_n383_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n471_), .B1(new_n474_), .B2(new_n403_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n467_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n461_), .B1(new_n453_), .B2(new_n448_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n447_), .A2(new_n448_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n445_), .B2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n402_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n460_), .A2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n452_), .A2(KEYINPUT33), .A3(new_n455_), .A4(new_n459_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n378_), .A2(KEYINPUT32), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n400_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n392_), .B2(new_n485_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n464_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n468_), .A2(new_n484_), .A3(new_n488_), .A4(new_n469_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n466_), .B1(new_n476_), .B2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G29gat), .B(G36gat), .Z(new_n491_));
  XOR2_X1   g290(.A(G43gat), .B(G50gat), .Z(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT15), .Z(new_n494_));
  XNOR2_X1  g293(.A(G1gat), .B(G8gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT72), .ZN(new_n496_));
  INV_X1    g295(.A(G22gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n407_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G15gat), .A2(G22gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G1gat), .A2(G8gat), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n498_), .A2(new_n499_), .B1(KEYINPUT14), .B2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n496_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n494_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n502_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n493_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n502_), .B(new_n493_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n503_), .A2(new_n508_), .B1(new_n509_), .B2(new_n505_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT75), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G169gat), .B(G197gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n510_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n490_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n521_));
  XOR2_X1   g320(.A(G71gat), .B(G78gat), .Z(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n521_), .A2(new_n522_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G85gat), .ZN(new_n526_));
  INV_X1    g325(.A(G92gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n530_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT8), .ZN(new_n538_));
  INV_X1    g337(.A(new_n536_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT9), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT65), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n529_), .A2(new_n541_), .A3(new_n540_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n529_), .B2(new_n540_), .ZN(new_n543_));
  OAI221_X1 g342(.A(new_n528_), .B1(new_n540_), .B2(new_n529_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT10), .B(G99gat), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT64), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n539_), .B(new_n544_), .C1(new_n547_), .C2(G106gat), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n525_), .B1(new_n538_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n518_), .B1(new_n549_), .B2(KEYINPUT12), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n537_), .A2(KEYINPUT8), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n537_), .A2(KEYINPUT8), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n545_), .B(KEYINPUT64), .ZN(new_n555_));
  INV_X1    g354(.A(G106gat), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n536_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n553_), .A2(new_n554_), .B1(new_n557_), .B2(new_n544_), .ZN(new_n558_));
  OAI211_X1 g357(.A(KEYINPUT66), .B(new_n551_), .C1(new_n558_), .C2(new_n525_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n550_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  INV_X1    g360(.A(new_n554_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n548_), .B1(new_n562_), .B2(new_n552_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n563_), .A2(KEYINPUT12), .A3(new_n524_), .A4(new_n523_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n558_), .A2(new_n525_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n565_), .ZN(new_n568_));
  OAI211_X1 g367(.A(G230gat), .B(G233gat), .C1(new_n568_), .C2(new_n549_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G120gat), .B(G148gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT5), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n574_), .B(KEYINPUT67), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n570_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n575_), .B1(new_n570_), .B2(new_n578_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n584_));
  INV_X1    g383(.A(new_n581_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n583_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT34), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT35), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT69), .Z(new_n591_));
  NAND3_X1  g390(.A1(new_n558_), .A2(KEYINPUT70), .A3(new_n507_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT70), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n563_), .B2(new_n493_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n589_), .A2(KEYINPUT35), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n494_), .B2(new_n563_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n591_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n595_), .A2(new_n597_), .A3(new_n591_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT36), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n599_), .A2(new_n600_), .A3(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n603_), .B(KEYINPUT36), .Z(new_n606_));
  INV_X1    g405(.A(new_n600_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n606_), .B1(new_n607_), .B2(new_n598_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n608_), .A3(KEYINPUT37), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(KEYINPUT71), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT71), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n612_), .B(new_n606_), .C1(new_n607_), .C2(new_n598_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n605_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n610_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n525_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n506_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT74), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT16), .ZN(new_n622_));
  XOR2_X1   g421(.A(G183gat), .B(G211gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n620_), .B1(new_n625_), .B2(KEYINPUT17), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n619_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(KEYINPUT73), .A3(KEYINPUT17), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(KEYINPUT17), .B2(new_n625_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n625_), .A2(KEYINPUT73), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n619_), .A2(new_n631_), .A3(new_n626_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n616_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n587_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n517_), .A2(KEYINPUT100), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT100), .B1(new_n517_), .B2(new_n635_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT101), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n636_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n471_), .A2(G1gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n639_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n639_), .A2(new_n642_), .A3(KEYINPUT38), .A4(new_n643_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n614_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n490_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n633_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n587_), .A2(new_n516_), .A3(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n471_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n646_), .A2(new_n647_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n646_), .A2(KEYINPUT102), .A3(new_n647_), .A4(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1324gat));
  INV_X1    g457(.A(G8gat), .ZN(new_n659_));
  INV_X1    g458(.A(new_n405_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n639_), .A2(new_n642_), .A3(new_n659_), .A4(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n652_), .A2(KEYINPUT103), .A3(new_n405_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n659_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT103), .B1(new_n652_), .B2(new_n405_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n664_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n661_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT40), .B(new_n661_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n652_), .B2(new_n437_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT41), .Z(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n637_), .A2(new_n638_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n407_), .A3(new_n467_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT105), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n675_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n676_), .A2(new_n679_), .A3(new_n680_), .ZN(G1326gat));
  OAI21_X1  g480(.A(G22gat), .B1(new_n652_), .B2(new_n293_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT42), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n677_), .A2(new_n497_), .A3(new_n470_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1327gat));
  NAND2_X1  g484(.A1(new_n648_), .A2(new_n650_), .ZN(new_n686_));
  NOR4_X1   g485(.A1(new_n490_), .A2(new_n516_), .A3(new_n587_), .A4(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(G29gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n464_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n490_), .B2(new_n616_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n293_), .A2(new_n405_), .A3(new_n465_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n464_), .B1(new_n399_), .B2(new_n404_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n437_), .B1(new_n697_), .B2(new_n293_), .ZN(new_n698_));
  AND4_X1   g497(.A1(new_n469_), .A2(new_n468_), .A3(new_n488_), .A4(new_n484_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n616_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n690_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n695_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n582_), .A2(new_n586_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n515_), .A3(new_n650_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n703_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  AOI211_X1 g507(.A(new_n708_), .B(new_n705_), .C1(new_n695_), .C2(new_n702_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n464_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G29gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n710_), .B2(new_n464_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n689_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  NAND2_X1  g514(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n716_));
  NOR2_X1   g515(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n687_), .A2(new_n718_), .A3(new_n660_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n719_), .A2(KEYINPUT45), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(KEYINPUT45), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT108), .B1(new_n710_), .B2(new_n660_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n489_), .B(new_n437_), .C1(new_n293_), .C2(new_n697_), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n616_), .B(new_n691_), .C1(new_n724_), .C2(new_n696_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n693_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n706_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n708_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT44), .B(new_n706_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n728_), .A2(KEYINPUT108), .A3(new_n660_), .A4(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G36gat), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n716_), .B(new_n722_), .C1(new_n723_), .C2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n728_), .A2(new_n660_), .A3(new_n729_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(G36gat), .A3(new_n730_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n716_), .B1(new_n737_), .B2(new_n722_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n733_), .A2(new_n738_), .ZN(G1329gat));
  NAND2_X1  g538(.A1(new_n710_), .A2(new_n467_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n437_), .A2(G43gat), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n740_), .A2(G43gat), .B1(new_n687_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n742_), .B(new_n744_), .ZN(G1330gat));
  AOI21_X1  g544(.A(G50gat), .B1(new_n687_), .B2(new_n470_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n470_), .A2(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n710_), .B2(new_n747_), .ZN(G1331gat));
  NOR4_X1   g547(.A1(new_n490_), .A2(new_n515_), .A3(new_n704_), .A4(new_n634_), .ZN(new_n749_));
  INV_X1    g548(.A(G57gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n464_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n704_), .A2(new_n515_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n649_), .A2(new_n633_), .A3(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT111), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(new_n464_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n755_), .B2(new_n750_), .ZN(G1332gat));
  INV_X1    g555(.A(G64gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n749_), .A2(new_n757_), .A3(new_n660_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(new_n660_), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(G64gat), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G64gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(G1333gat));
  INV_X1    g562(.A(G71gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n749_), .A2(new_n764_), .A3(new_n467_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n754_), .A2(new_n467_), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(G71gat), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G71gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(G1334gat));
  NOR2_X1   g569(.A1(new_n293_), .A2(G78gat), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT114), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n749_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n754_), .A2(new_n470_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G78gat), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(KEYINPUT50), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(KEYINPUT50), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(G1335gat));
  NOR3_X1   g577(.A1(new_n704_), .A2(new_n515_), .A3(new_n633_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n703_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780_), .B2(new_n471_), .ZN(new_n781_));
  NOR4_X1   g580(.A1(new_n490_), .A2(new_n515_), .A3(new_n704_), .A4(new_n686_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n526_), .A3(new_n464_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n780_), .B2(new_n405_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n527_), .A3(new_n660_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1337gat));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n703_), .A2(new_n467_), .A3(new_n779_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n437_), .A2(new_n547_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n789_), .A2(G99gat), .B1(new_n782_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT51), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n791_), .B2(new_n788_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n794_), .B1(new_n793_), .B2(new_n796_), .ZN(G1338gat));
  NAND3_X1  g596(.A1(new_n782_), .A2(new_n556_), .A3(new_n470_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n703_), .A2(new_n470_), .A3(new_n779_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  AND4_X1   g600(.A1(new_n799_), .A2(new_n800_), .A3(new_n801_), .A4(G106gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n556_), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n800_), .A2(new_n803_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n798_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g605(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n635_), .A2(new_n516_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n807_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n704_), .A2(new_n633_), .A3(new_n616_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n515_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n561_), .B1(new_n560_), .B2(new_n566_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n567_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n560_), .A2(new_n566_), .A3(KEYINPUT55), .A4(new_n561_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n577_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n820_), .B(new_n578_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n515_), .B(new_n575_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n510_), .A2(new_n514_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n503_), .B(new_n505_), .C1(new_n502_), .C2(new_n493_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n514_), .B1(new_n509_), .B2(new_n504_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n583_), .A2(new_n823_), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n648_), .B1(new_n822_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n813_), .B1(new_n828_), .B2(KEYINPUT57), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n575_), .A2(new_n515_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n818_), .A2(new_n577_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n820_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n830_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n827_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n614_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(KEYINPUT119), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n828_), .A2(KEYINPUT57), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n575_), .A2(new_n823_), .A3(new_n826_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n840_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n616_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n832_), .A2(new_n833_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n841_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n845_), .A3(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n829_), .A2(new_n838_), .A3(new_n839_), .A4(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n812_), .B1(new_n849_), .B2(new_n650_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n293_), .A2(new_n405_), .A3(new_n464_), .A4(new_n467_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(G113gat), .B1(new_n852_), .B2(new_n515_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n836_), .A2(new_n837_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n848_), .A2(new_n854_), .A3(new_n839_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(KEYINPUT121), .A3(new_n650_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT121), .B1(new_n855_), .B2(new_n650_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n812_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n851_), .A2(KEYINPUT59), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n852_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n516_), .A2(KEYINPUT122), .ZN(new_n866_));
  MUX2_X1   g665(.A(KEYINPUT122), .B(new_n866_), .S(G113gat), .Z(new_n867_));
  AOI21_X1  g666(.A(new_n853_), .B1(new_n865_), .B2(new_n867_), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n704_), .B2(KEYINPUT60), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(KEYINPUT60), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(KEYINPUT123), .B2(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n852_), .B(new_n872_), .C1(KEYINPUT123), .C2(new_n870_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n862_), .A2(new_n864_), .A3(new_n704_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n869_), .ZN(G1341gat));
  OAI21_X1  g674(.A(KEYINPUT59), .B1(new_n850_), .B2(new_n851_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(new_n633_), .C1(new_n859_), .C2(new_n861_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G127gat), .ZN(new_n878_));
  INV_X1    g677(.A(G127gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n852_), .A2(new_n879_), .A3(new_n633_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT124), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n878_), .A2(new_n883_), .A3(new_n880_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1342gat));
  INV_X1    g684(.A(G134gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n852_), .A2(new_n886_), .A3(new_n648_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n862_), .A2(new_n864_), .A3(new_n616_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n886_), .ZN(G1343gat));
  NOR3_X1   g688(.A1(new_n850_), .A2(new_n293_), .A3(new_n467_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n660_), .A2(new_n471_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n516_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n704_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g695(.A1(new_n892_), .A2(new_n650_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  XOR2_X1   g697(.A(new_n897_), .B(new_n898_), .Z(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n892_), .B2(new_n616_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n614_), .A2(G162gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n892_), .B2(new_n901_), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n405_), .A2(new_n464_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n467_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n859_), .A2(new_n470_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n515_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n906_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  NOR4_X1   g707(.A1(new_n859_), .A2(new_n470_), .A3(new_n516_), .A4(new_n904_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n296_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n907_), .B(new_n910_), .C1(new_n360_), .C2(new_n906_), .ZN(G1348gat));
  AOI21_X1  g710(.A(G176gat), .B1(new_n905_), .B2(new_n587_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n850_), .A2(new_n470_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n904_), .A2(new_n297_), .A3(new_n704_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1349gat));
  NOR2_X1   g714(.A1(new_n650_), .A2(new_n352_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n913_), .A2(new_n467_), .A3(new_n633_), .A4(new_n903_), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n905_), .A2(new_n916_), .B1(new_n917_), .B2(new_n324_), .ZN(G1350gat));
  NAND4_X1  g717(.A1(new_n905_), .A2(new_n351_), .A3(new_n353_), .A4(new_n648_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n905_), .A2(new_n701_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n310_), .ZN(G1351gat));
  INV_X1    g720(.A(new_n903_), .ZN(new_n922_));
  NOR4_X1   g721(.A1(new_n850_), .A2(new_n293_), .A3(new_n467_), .A4(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n515_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g724(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT125), .B(G204gat), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n923_), .A2(new_n587_), .ZN(new_n928_));
  MUX2_X1   g727(.A(new_n926_), .B(new_n927_), .S(new_n928_), .Z(G1353gat));
  NAND2_X1  g728(.A1(new_n923_), .A2(new_n633_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  AND2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n933_), .B1(new_n930_), .B2(new_n931_), .ZN(G1354gat));
  NAND2_X1  g733(.A1(new_n923_), .A2(new_n648_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT126), .B(G218gat), .Z(new_n936_));
  NOR2_X1   g735(.A1(new_n616_), .A2(new_n936_), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n935_), .A2(new_n936_), .B1(new_n923_), .B2(new_n937_), .ZN(G1355gat));
endmodule


