//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207_));
  INV_X1    g006(.A(G134gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G127gat), .ZN(new_n209_));
  INV_X1    g008(.A(G127gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G134gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G120gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G113gat), .ZN(new_n214_));
  INV_X1    g013(.A(G113gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G120gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n209_), .A2(new_n211_), .A3(new_n214_), .A4(new_n216_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G141gat), .B(G148gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT89), .A2(G155gat), .A3(G162gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT1), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G155gat), .A3(G162gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n222_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233_));
  INV_X1    g032(.A(G141gat), .ZN(new_n234_));
  INV_X1    g033(.A(G148gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G141gat), .A2(G148gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n236_), .A2(new_n239_), .A3(new_n240_), .A4(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n227_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT89), .ZN(new_n244_));
  INV_X1    g043(.A(G155gat), .ZN(new_n245_));
  INV_X1    g044(.A(G162gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n247_), .B2(new_n223_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n242_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n220_), .B1(new_n232_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n207_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n218_), .A2(new_n219_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n242_), .A2(new_n248_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n228_), .A2(new_n230_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n247_), .A2(new_n223_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n221_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n253_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n232_), .A2(new_n249_), .A3(new_n220_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT4), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT99), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n252_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(new_n259_), .A3(new_n207_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n261_), .B1(new_n252_), .B2(new_n260_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n206_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n258_), .A2(KEYINPUT4), .A3(new_n259_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n207_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(new_n258_), .B2(KEYINPUT4), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT99), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n206_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n263_), .A4(new_n262_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(G15gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT30), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT31), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT23), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT87), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT23), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n280_), .B(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n284_), .B2(KEYINPUT87), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(G183gat), .B2(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT22), .B(G169gat), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT86), .ZN(new_n290_));
  INV_X1    g089(.A(G169gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT22), .ZN(new_n292_));
  AOI21_X1  g091(.A(G176gat), .B1(new_n292_), .B2(KEYINPUT86), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n288_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n286_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G176gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n287_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(KEYINPUT24), .B2(new_n297_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(new_n284_), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT84), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G190gat), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n302_), .A2(new_n303_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n305_), .A2(G190gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n309_), .B(new_n310_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n300_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n295_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G71gat), .B(G99gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT88), .B(G43gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n313_), .A2(new_n316_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n253_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n318_), .A2(new_n253_), .A3(new_n319_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n279_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n322_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(new_n278_), .A3(new_n320_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n273_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT21), .B1(new_n327_), .B2(KEYINPUT95), .ZN(new_n328_));
  INV_X1    g127(.A(G218gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G211gat), .ZN(new_n330_));
  INV_X1    g129(.A(G211gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G218gat), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n330_), .A2(new_n332_), .A3(KEYINPUT95), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT92), .ZN(new_n335_));
  INV_X1    g134(.A(G204gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(G197gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(G197gat), .ZN(new_n338_));
  INV_X1    g137(.A(G197gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n338_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT21), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n327_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n344_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n330_), .A2(new_n332_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n339_), .A2(G204gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n338_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(KEYINPUT21), .B2(new_n352_), .ZN(new_n353_));
  AND2_X1   g152(.A1(KEYINPUT93), .A2(KEYINPUT21), .ZN(new_n354_));
  NOR2_X1   g153(.A1(KEYINPUT93), .A2(KEYINPUT21), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n356_), .A2(new_n337_), .A3(new_n338_), .A4(new_n340_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT94), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n342_), .B1(new_n349_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT96), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n348_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n353_), .A2(KEYINPUT94), .A3(new_n357_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n361_), .A2(new_n362_), .B1(new_n341_), .B2(new_n334_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT96), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT91), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n232_), .A2(new_n249_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(KEYINPUT29), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n360_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n368_), .A2(KEYINPUT29), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n367_), .B1(new_n363_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT97), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n368_), .A2(KEYINPUT29), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n377_), .B(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n370_), .A2(new_n374_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n371_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n375_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n376_), .A2(new_n384_), .A3(new_n375_), .A4(new_n381_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n295_), .A2(new_n312_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n360_), .A2(new_n365_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n399_));
  AND4_X1   g198(.A1(new_n302_), .A2(new_n309_), .A3(new_n310_), .A4(new_n306_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(new_n299_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n284_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(G183gat), .B2(G190gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n288_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n401_), .A2(new_n285_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n399_), .B1(new_n363_), .B2(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n395_), .A2(new_n398_), .A3(new_n406_), .ZN(new_n407_));
  AOI221_X4 g206(.A(KEYINPUT96), .B1(new_n334_), .B2(new_n341_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n361_), .A2(new_n362_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n364_), .B1(new_n409_), .B2(new_n342_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n313_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n405_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n399_), .B1(new_n412_), .B2(new_n359_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n398_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n393_), .B1(new_n407_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n394_), .B1(new_n360_), .B2(new_n365_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT20), .B1(new_n363_), .B2(new_n405_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n397_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n395_), .A2(new_n398_), .A3(new_n406_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n393_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n415_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT27), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n416_), .A2(new_n397_), .A3(new_n417_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n398_), .B1(new_n395_), .B2(new_n406_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n393_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(KEYINPUT27), .A3(new_n421_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n326_), .A2(new_n388_), .A3(new_n424_), .A4(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT104), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n323_), .A2(new_n325_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n387_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n376_), .A2(new_n381_), .B1(new_n384_), .B2(new_n375_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n273_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n424_), .A4(new_n428_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT101), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n268_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n440_), .A2(new_n260_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n258_), .A2(new_n259_), .A3(new_n268_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n206_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n439_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n260_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n445_), .A2(KEYINPUT101), .A3(new_n206_), .A4(new_n442_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n272_), .A2(new_n438_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n264_), .A2(new_n265_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(KEYINPUT33), .A3(new_n271_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n415_), .A2(new_n421_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n420_), .A2(KEYINPUT32), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n418_), .A2(new_n419_), .A3(new_n451_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n273_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT102), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n388_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n437_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n456_), .B2(new_n388_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n432_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT103), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT103), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n463_), .B(new_n432_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n430_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G29gat), .B(G36gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G43gat), .B(G50gat), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n467_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473_));
  INV_X1    g272(.A(G1gat), .ZN(new_n474_));
  INV_X1    g273(.A(G8gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G8gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n472_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n479_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n470_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(new_n469_), .A3(new_n468_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(KEYINPUT82), .A3(new_n485_), .ZN(new_n486_));
  OR3_X1    g285(.A1(new_n482_), .A2(KEYINPUT82), .A3(new_n470_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n481_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n486_), .A2(new_n487_), .A3(KEYINPUT83), .A4(new_n488_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n484_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G113gat), .B(G141gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G169gat), .B(G197gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n493_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n465_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G85gat), .ZN(new_n500_));
  INV_X1    g299(.A(G92gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n504_), .B(new_n505_), .C1(new_n508_), .C2(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n502_), .A2(new_n503_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n506_), .B(KEYINPUT7), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n509_), .B(KEYINPUT6), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n513_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n512_), .B(KEYINPUT68), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT65), .ZN(new_n520_));
  AND3_X1   g319(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT66), .B1(new_n521_), .B2(new_n503_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n520_), .B(new_n522_), .C1(KEYINPUT66), .C2(new_n521_), .ZN(new_n523_));
  INV_X1    g322(.A(G106gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT64), .ZN(new_n526_));
  NAND2_X1  g325(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n524_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n523_), .A2(new_n515_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT68), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n516_), .A2(new_n532_), .A3(new_n505_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n518_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT69), .B(G71gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G78gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n536_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G78gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n535_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n538_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n534_), .A2(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n546_), .A2(KEYINPUT12), .ZN(new_n547_));
  INV_X1    g346(.A(new_n545_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n548_), .A2(new_n518_), .A3(new_n533_), .A4(new_n531_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT12), .A3(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n546_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT5), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT70), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n563_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT72), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n534_), .A2(new_n472_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT74), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n534_), .A2(new_n472_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(KEYINPUT35), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n518_), .A2(new_n531_), .A3(new_n470_), .A4(new_n533_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n574_), .A2(new_n576_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(KEYINPUT35), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n582_), .B(KEYINPUT76), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n573_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n580_), .A2(new_n579_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G190gat), .B(G218gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n591_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT36), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT75), .Z(new_n595_));
  NAND3_X1  g394(.A1(new_n584_), .A2(new_n589_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT77), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n588_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n592_), .A2(new_n593_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT36), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT78), .B1(new_n599_), .B2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n599_), .A2(KEYINPUT77), .A3(new_n595_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT78), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n587_), .B1(KEYINPUT74), .B2(new_n573_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n582_), .B1(new_n606_), .B2(new_n576_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n605_), .B(new_n601_), .C1(new_n607_), .C2(new_n588_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n598_), .A2(new_n603_), .A3(new_n604_), .A4(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT37), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT79), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n601_), .B1(new_n607_), .B2(new_n588_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(new_n596_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n610_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n611_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G183gat), .B(G211gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT17), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(KEYINPUT81), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n479_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n625_), .A2(KEYINPUT81), .A3(new_n482_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(G231gat), .A3(G233gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n631_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n545_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n623_), .A2(new_n624_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n548_), .A3(new_n632_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n618_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n572_), .A2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n499_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n474_), .A3(new_n273_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT38), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n613_), .B(KEYINPUT105), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n465_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n571_), .A2(new_n498_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n637_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n436_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n641_), .A2(new_n642_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n643_), .A2(new_n648_), .A3(new_n649_), .ZN(G1324gat));
  NAND2_X1  g449(.A1(new_n424_), .A2(new_n428_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n499_), .A2(new_n475_), .A3(new_n651_), .A4(new_n639_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT106), .Z(new_n653_));
  INV_X1    g452(.A(new_n651_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G8gat), .B1(new_n647_), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n656_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n653_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n653_), .A2(new_n657_), .A3(KEYINPUT40), .A4(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n647_), .B2(new_n432_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  NAND3_X1  g464(.A1(new_n640_), .A2(new_n275_), .A3(new_n431_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1326gat));
  OAI21_X1  g466(.A(G22gat), .B1(new_n647_), .B2(new_n388_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT42), .ZN(new_n669_));
  INV_X1    g468(.A(G22gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n640_), .A2(new_n670_), .A3(new_n435_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(new_n637_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n613_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n571_), .A2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n499_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n273_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n610_), .A2(new_n615_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT79), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n610_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n678_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n684_), .B1(new_n465_), .B2(new_n618_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n430_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n464_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n456_), .A2(new_n388_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT102), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n437_), .A3(new_n458_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n463_), .B1(new_n690_), .B2(new_n432_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n686_), .B1(new_n687_), .B2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n683_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT43), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n682_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n685_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n646_), .A2(new_n673_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT44), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n700_), .B(new_n697_), .C1(new_n685_), .C2(new_n695_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n273_), .A2(G29gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n677_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n702_), .B2(new_n651_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n499_), .A2(new_n706_), .A3(new_n651_), .A4(new_n675_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT45), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n707_), .B2(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n699_), .A2(new_n701_), .A3(new_n654_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT46), .B(new_n709_), .C1(new_n712_), .C2(new_n706_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1329gat));
  NAND3_X1  g513(.A1(new_n499_), .A2(new_n431_), .A3(new_n675_), .ZN(new_n715_));
  INV_X1    g514(.A(G43gat), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n696_), .A2(new_n698_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n700_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n696_), .A2(KEYINPUT44), .A3(new_n698_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n721_), .A2(G43gat), .A3(new_n431_), .A4(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n719_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n719_), .B2(new_n723_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n676_), .B2(new_n435_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n435_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n702_), .B2(new_n729_), .ZN(G1331gat));
  AND2_X1   g529(.A1(new_n637_), .A2(new_n498_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n645_), .A2(new_n572_), .A3(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT112), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(G57gat), .A3(new_n273_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n733_), .A2(KEYINPUT113), .A3(G57gat), .A4(new_n273_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  INV_X1    g537(.A(new_n570_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n567_), .ZN(new_n740_));
  NOR4_X1   g539(.A1(new_n465_), .A2(new_n638_), .A3(new_n497_), .A4(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n273_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n738_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n736_), .A2(new_n737_), .A3(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(G64gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n741_), .A2(new_n747_), .A3(new_n651_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n733_), .A2(new_n651_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G64gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT48), .B(new_n747_), .C1(new_n733_), .C2(new_n651_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1333gat));
  INV_X1    g552(.A(G71gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n741_), .A2(new_n754_), .A3(new_n431_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n645_), .A2(new_n572_), .A3(new_n731_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(KEYINPUT112), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT112), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n431_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n756_), .B1(new_n760_), .B2(G71gat), .ZN(new_n761_));
  AOI211_X1 g560(.A(KEYINPUT49), .B(new_n754_), .C1(new_n733_), .C2(new_n431_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n755_), .B1(new_n761_), .B2(new_n762_), .ZN(G1334gat));
  NAND3_X1  g562(.A1(new_n741_), .A2(new_n541_), .A3(new_n435_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n733_), .A2(new_n435_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G78gat), .ZN(new_n767_));
  AOI211_X1 g566(.A(KEYINPUT50), .B(new_n541_), .C1(new_n733_), .C2(new_n435_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(G1335gat));
  NOR3_X1   g568(.A1(new_n740_), .A2(new_n497_), .A3(new_n637_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n696_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(G85gat), .A3(new_n273_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n572_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n674_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n465_), .A2(new_n497_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n500_), .B1(new_n776_), .B2(new_n436_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT114), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(KEYINPUT114), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n772_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n772_), .B(KEYINPUT115), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1336gat));
  INV_X1    g583(.A(new_n776_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n501_), .A3(new_n651_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n771_), .A2(new_n651_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n501_), .ZN(G1337gat));
  OAI21_X1  g587(.A(new_n431_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n776_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n771_), .A2(new_n431_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G99gat), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT51), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n792_), .B(new_n794_), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n785_), .A2(new_n524_), .A3(new_n435_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n696_), .A2(new_n435_), .A3(new_n770_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G106gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n796_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  XOR2_X1   g604(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n547_), .A2(new_n550_), .A3(new_n555_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n553_), .A2(KEYINPUT55), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n555_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n562_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n809_), .A2(KEYINPUT56), .A3(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n486_), .A2(new_n487_), .A3(new_n481_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n481_), .B1(new_n482_), .B2(new_n470_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n496_), .B1(new_n480_), .B2(new_n819_), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n493_), .A2(new_n496_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n553_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n817_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n817_), .A2(KEYINPUT58), .A3(new_n823_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n826_), .B(new_n827_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n613_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n809_), .A2(new_n812_), .A3(KEYINPUT117), .A4(KEYINPUT56), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n830_), .A2(new_n497_), .A3(new_n822_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n815_), .A2(new_n832_), .A3(new_n816_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n564_), .A2(new_n565_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n835_), .A2(new_n821_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT57), .B(new_n829_), .C1(new_n834_), .C2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n831_), .A2(new_n833_), .B1(new_n835_), .B2(new_n821_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n613_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n828_), .A2(new_n837_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n618_), .A2(new_n842_), .A3(new_n740_), .A4(new_n731_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n740_), .A2(new_n731_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT54), .B1(new_n682_), .B2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n673_), .A2(new_n841_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n651_), .A2(new_n435_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n431_), .A3(new_n273_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n807_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n841_), .A2(new_n673_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n843_), .A2(new_n845_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n848_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n849_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT119), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n849_), .A2(new_n855_), .A3(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n497_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G113gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n852_), .A2(new_n853_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n215_), .A3(new_n497_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n864_), .ZN(G1340gat));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n856_), .B2(new_n773_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n740_), .B2(G120gat), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n863_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n849_), .A2(new_n855_), .A3(KEYINPUT120), .A4(new_n572_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G120gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n863_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1341gat));
  OAI21_X1  g674(.A(new_n210_), .B1(new_n862_), .B2(new_n673_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT121), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n857_), .A2(new_n859_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n637_), .A2(G127gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT122), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n877_), .B1(new_n878_), .B2(new_n880_), .ZN(G1342gat));
  NAND3_X1  g680(.A1(new_n857_), .A2(new_n682_), .A3(new_n859_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G134gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n863_), .A2(new_n208_), .A3(new_n644_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1343gat));
  NOR3_X1   g684(.A1(new_n431_), .A2(new_n388_), .A3(new_n436_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n852_), .A2(new_n654_), .A3(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n498_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n234_), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n773_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n235_), .ZN(G1345gat));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n673_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT61), .B(G155gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  INV_X1    g693(.A(new_n644_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n246_), .B1(new_n887_), .B2(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT123), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n887_), .A2(new_n246_), .A3(new_n618_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1347gat));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n852_), .A2(new_n388_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n651_), .A2(new_n326_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT124), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n498_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n900_), .B1(new_n906_), .B2(new_n291_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n289_), .ZN(new_n908_));
  OAI211_X1 g707(.A(KEYINPUT62), .B(G169gat), .C1(new_n905_), .C2(new_n498_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n904_), .B2(new_n571_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n901_), .B(KEYINPUT125), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n773_), .A2(new_n296_), .A3(new_n903_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT126), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n912_), .A2(new_n916_), .A3(new_n913_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n911_), .B1(new_n915_), .B2(new_n917_), .ZN(G1349gat));
  NAND2_X1  g717(.A1(new_n302_), .A2(new_n310_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n904_), .A2(new_n919_), .A3(new_n637_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n903_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n912_), .A2(new_n637_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n922_), .B2(new_n301_), .ZN(G1350gat));
  OAI21_X1  g722(.A(G190gat), .B1(new_n905_), .B2(new_n618_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n644_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n905_), .B2(new_n925_), .ZN(G1351gat));
  NAND3_X1  g725(.A1(new_n435_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n846_), .A2(new_n654_), .A3(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n497_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n572_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g731(.A1(new_n928_), .A2(new_n637_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  AND2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n936_), .B1(new_n933_), .B2(new_n934_), .ZN(G1354gat));
  NAND2_X1  g736(.A1(new_n928_), .A2(new_n644_), .ZN(new_n938_));
  XOR2_X1   g737(.A(KEYINPUT127), .B(G218gat), .Z(new_n939_));
  NOR2_X1   g738(.A1(new_n618_), .A2(new_n939_), .ZN(new_n940_));
  AOI22_X1  g739(.A1(new_n938_), .A2(new_n939_), .B1(new_n928_), .B2(new_n940_), .ZN(G1355gat));
endmodule


