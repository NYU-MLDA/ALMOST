//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_;
  INV_X1    g000(.A(G155gat), .ZN(new_n202_));
  INV_X1    g001(.A(G162gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT83), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(G155gat), .B2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n211_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n208_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT84), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n208_), .A2(new_n217_), .A3(KEYINPUT84), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT82), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n212_), .B1(new_n209_), .B2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n224_), .B1(new_n223_), .B2(new_n209_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n207_), .B(KEYINPUT1), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n204_), .A2(new_n206_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n222_), .A2(KEYINPUT85), .A3(new_n228_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT28), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT28), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(new_n237_), .A3(new_n234_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G22gat), .B(G50gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n239_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n237_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n242_));
  AOI211_X1 g041(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n231_), .C2(new_n232_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT90), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G211gat), .B(G218gat), .Z(new_n248_));
  INV_X1    g047(.A(KEYINPUT21), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G197gat), .B(G204gat), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G197gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(G197gat), .B(G204gat), .Z(new_n254_));
  OAI211_X1 g053(.A(KEYINPUT21), .B(new_n253_), .C1(new_n254_), .C2(KEYINPUT87), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT88), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT88), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n255_), .A3(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n250_), .A2(new_n249_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n257_), .A2(new_n259_), .B1(new_n248_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(KEYINPUT29), .B2(new_n229_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G228gat), .A2(G233gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT89), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n229_), .A2(KEYINPUT29), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT89), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(G228gat), .A4(G233gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT86), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT86), .A4(KEYINPUT29), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n265_), .A4(new_n263_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G78gat), .B(G106gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n240_), .A2(new_n244_), .A3(KEYINPUT90), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n270_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n247_), .A2(new_n278_), .A3(new_n279_), .A4(new_n280_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n270_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n276_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n246_), .B(new_n245_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G127gat), .B(G134gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n231_), .A2(new_n232_), .A3(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n229_), .A2(new_n288_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT4), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT4), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n293_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G1gat), .B(G29gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G57gat), .B(G85gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n299_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT27), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT23), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(G183gat), .B2(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT77), .B(G176gat), .ZN(new_n315_));
  INV_X1    g114(.A(G169gat), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT22), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(KEYINPUT22), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT76), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n313_), .B(new_n314_), .C1(new_n318_), .C2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n322_), .A2(KEYINPUT75), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(KEYINPUT75), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT24), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT25), .B(G183gat), .ZN(new_n328_));
  INV_X1    g127(.A(G190gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT26), .B1(new_n329_), .B2(KEYINPUT74), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(KEYINPUT26), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n328_), .B(new_n330_), .C1(new_n331_), .C2(KEYINPUT74), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n323_), .A2(KEYINPUT24), .A3(new_n324_), .A4(new_n314_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n327_), .A2(new_n332_), .A3(new_n312_), .A4(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n321_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT78), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n321_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n261_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(KEYINPUT26), .B(G190gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT92), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n328_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n322_), .A2(new_n326_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n333_), .A2(new_n312_), .A3(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n314_), .B(KEYINPUT93), .Z(new_n345_));
  AND2_X1   g144(.A1(new_n317_), .A2(new_n319_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n315_), .B2(new_n346_), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n342_), .A2(new_n344_), .B1(new_n313_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT20), .B1(new_n261_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n310_), .B1(new_n339_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n336_), .A2(new_n338_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n265_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n310_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n261_), .B2(new_n348_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT18), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  AND3_X1   g159(.A1(new_n350_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n350_), .B2(new_n356_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n307_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n360_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n339_), .A2(new_n349_), .A3(new_n310_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n353_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n350_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(KEYINPUT27), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n297_), .A2(new_n304_), .A3(new_n298_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n306_), .A2(new_n363_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT96), .B1(new_n285_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT96), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n284_), .A4(new_n281_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n362_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n294_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n304_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n376_), .B(new_n368_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n304_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(KEYINPUT95), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n381_), .B2(KEYINPUT33), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n380_), .A2(KEYINPUT95), .A3(KEYINPUT33), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n306_), .A2(new_n370_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n365_), .A2(new_n366_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(KEYINPUT32), .A3(new_n360_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n350_), .A2(new_n356_), .A3(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n382_), .A2(new_n383_), .B1(new_n384_), .B2(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n281_), .A2(new_n284_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n372_), .B(new_n375_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393_));
  INV_X1    g192(.A(G43gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(G15gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n395_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n351_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n399_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n351_), .B(KEYINPUT30), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT79), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n403_), .A2(new_n405_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n288_), .B(KEYINPUT81), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT80), .B1(new_n408_), .B2(KEYINPUT31), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n409_), .B1(KEYINPUT31), .B2(new_n408_), .ZN(new_n410_));
  OR3_X1    g209(.A1(new_n406_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n363_), .A2(new_n369_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT97), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n413_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI211_X1 g217(.A(KEYINPUT97), .B(new_n415_), .C1(new_n281_), .C2(new_n284_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n384_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n392_), .A2(new_n414_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G113gat), .B(G141gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G169gat), .B(G197gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G29gat), .B(G36gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT70), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G43gat), .B(G50gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n427_), .A2(KEYINPUT70), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(KEYINPUT70), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n429_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G15gat), .B(G22gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT71), .B(G8gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G1gat), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n439_), .B2(KEYINPUT14), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT72), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G8gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n440_), .B(KEYINPUT72), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(new_n443_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n436_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n443_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n444_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n431_), .A2(KEYINPUT15), .A3(new_n434_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT15), .B1(new_n431_), .B2(new_n434_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n450_), .B(new_n451_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n448_), .A2(new_n449_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n451_), .A3(new_n435_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n449_), .B1(new_n448_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n426_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n448_), .A2(new_n449_), .A3(new_n454_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n450_), .A2(new_n451_), .A3(new_n435_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n435_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n459_), .B(new_n425_), .C1(new_n462_), .C2(new_n449_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT73), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(KEYINPUT73), .B(new_n426_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n422_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G230gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT64), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G99gat), .A2(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G85gat), .ZN(new_n481_));
  INV_X1    g280(.A(G92gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(KEYINPUT9), .A3(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(KEYINPUT9), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n476_), .A2(new_n480_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT8), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(G99gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n478_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n474_), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n490_), .B(new_n493_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n483_), .A2(new_n484_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n489_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n489_), .A3(new_n498_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n488_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G71gat), .B(G78gat), .ZN(new_n503_));
  INV_X1    g302(.A(G64gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G57gat), .ZN(new_n505_));
  INV_X1    g304(.A(G57gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G64gat), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n503_), .A2(KEYINPUT11), .A3(new_n505_), .A4(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n507_), .A3(KEYINPUT11), .ZN(new_n509_));
  INV_X1    g308(.A(G78gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(G71gat), .ZN(new_n511_));
  INV_X1    g310(.A(G71gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G78gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n509_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT11), .B1(new_n505_), .B2(new_n507_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n508_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT65), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT65), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n508_), .B(new_n519_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n502_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n471_), .B1(new_n522_), .B2(KEYINPUT66), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(KEYINPUT66), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n502_), .A2(new_n521_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n520_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n505_), .A2(new_n507_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT11), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(new_n509_), .A3(new_n514_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n519_), .B1(new_n532_), .B2(new_n508_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n490_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AOI211_X1 g336(.A(KEYINPUT8), .B(new_n497_), .C1(new_n537_), .C2(new_n476_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n487_), .B1(new_n538_), .B2(new_n499_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n471_), .B1(new_n534_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT68), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT68), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n525_), .A2(new_n542_), .A3(new_n471_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT67), .B(new_n487_), .C1(new_n538_), .C2(new_n499_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n532_), .A2(KEYINPUT12), .A3(new_n508_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n502_), .B2(new_n521_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n544_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G120gat), .B(G148gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n527_), .A2(new_n554_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n559_), .B1(new_n527_), .B2(new_n554_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT13), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(KEYINPUT13), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n450_), .A2(new_n451_), .ZN(new_n568_));
  AND2_X1   g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(new_n517_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572_));
  XOR2_X1   g371(.A(G127gat), .B(G155gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n571_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n570_), .B2(new_n517_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n576_), .B(new_n572_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n570_), .B2(new_n534_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n570_), .B2(new_n534_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n436_), .A2(new_n502_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n546_), .A2(new_n547_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n452_), .A2(new_n453_), .ZN(new_n588_));
  OAI221_X1 g387(.A(new_n584_), .B1(KEYINPUT35), .B2(new_n586_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n594_), .B(KEYINPUT36), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n591_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT37), .B1(new_n597_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n596_), .B(new_n602_), .C1(new_n591_), .C2(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n583_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n567_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n468_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(G1gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n384_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n607_), .A2(KEYINPUT98), .A3(new_n608_), .A4(new_n384_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(KEYINPUT38), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT99), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n597_), .A2(new_n600_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n375_), .A2(new_n372_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT33), .B1(new_n380_), .B2(KEYINPUT95), .ZN(new_n617_));
  INV_X1    g416(.A(new_n379_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n383_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n389_), .A2(new_n384_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n391_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n414_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT97), .B1(new_n391_), .B2(new_n415_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n416_), .A2(new_n417_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n623_), .A2(new_n421_), .A3(new_n624_), .A4(new_n413_), .ZN(new_n625_));
  AOI211_X1 g424(.A(new_n582_), .B(new_n615_), .C1(new_n622_), .C2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n567_), .A2(new_n467_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT100), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n421_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n611_), .A2(new_n612_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT101), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n632_), .A2(KEYINPUT101), .A3(new_n633_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n614_), .B(new_n631_), .C1(new_n634_), .C2(new_n635_), .ZN(G1324gat));
  NAND2_X1  g435(.A1(new_n628_), .A2(new_n415_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n637_), .B2(G8gat), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n415_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n438_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n607_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n642_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n642_), .B2(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1325gat));
  AOI21_X1  g450(.A(new_n397_), .B1(new_n629_), .B2(new_n413_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT41), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n607_), .A2(new_n397_), .A3(new_n413_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1326gat));
  INV_X1    g454(.A(G22gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n285_), .B(KEYINPUT103), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n629_), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n607_), .A2(new_n656_), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1327gat));
  NAND2_X1  g462(.A1(new_n582_), .A2(new_n615_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n567_), .A2(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n468_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n384_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n627_), .A2(new_n582_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n669_), .B(KEYINPUT43), .C1(new_n422_), .C2(new_n604_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n604_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(KEYINPUT105), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n668_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT44), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n384_), .A2(G29gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n667_), .B1(new_n678_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  OAI21_X1  g480(.A(G36gat), .B1(new_n677_), .B2(new_n644_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(G36gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n666_), .A2(new_n684_), .A3(new_n415_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT45), .Z(new_n686_));
  OAI21_X1  g485(.A(new_n681_), .B1(new_n683_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n686_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(KEYINPUT46), .A3(new_n682_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1329gat));
  NAND3_X1  g489(.A1(new_n678_), .A2(G43gat), .A3(new_n413_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n666_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n394_), .B1(new_n692_), .B2(new_n414_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n691_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n666_), .B2(new_n658_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n391_), .A2(G50gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n678_), .B2(new_n699_), .ZN(G1331gat));
  INV_X1    g499(.A(new_n467_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n566_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n626_), .A2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT108), .ZN(new_n704_));
  OAI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n421_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n422_), .A2(new_n701_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n706_), .A2(new_n583_), .A3(new_n604_), .A4(new_n567_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n506_), .A3(new_n384_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(G1332gat));
  OAI21_X1  g509(.A(G64gat), .B1(new_n704_), .B2(new_n644_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(new_n504_), .A3(new_n415_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n704_), .B2(new_n414_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n708_), .A2(new_n512_), .A3(new_n413_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n704_), .B2(new_n657_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n708_), .A2(new_n510_), .A3(new_n658_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1335gat));
  NAND2_X1  g521(.A1(new_n702_), .A2(new_n582_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n421_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n706_), .A2(new_n582_), .A3(new_n615_), .A4(new_n567_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(new_n481_), .A3(new_n384_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT109), .ZN(G1336gat));
  OAI21_X1  g530(.A(G92gat), .B1(new_n725_), .B2(new_n644_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n728_), .A2(new_n482_), .A3(new_n415_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n725_), .B2(new_n414_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n413_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n727_), .B2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g537(.A1(new_n728_), .A2(new_n478_), .A3(new_n391_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  AOI211_X1 g539(.A(new_n285_), .B(new_n723_), .C1(new_n670_), .C2(new_n673_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n478_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n724_), .B2(new_n391_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n740_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n670_), .A2(new_n673_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n723_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n747_), .A2(new_n742_), .A3(new_n391_), .A4(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G106gat), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n750_), .A2(new_n744_), .A3(KEYINPUT52), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n739_), .B1(new_n746_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(new_n739_), .C1(new_n746_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  NAND2_X1  g555(.A1(new_n606_), .A2(new_n467_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n559_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n544_), .A2(new_n553_), .A3(KEYINPUT55), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n550_), .A2(new_n552_), .A3(new_n525_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n470_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT55), .B1(new_n544_), .B2(new_n553_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n761_), .B(new_n763_), .C1(new_n764_), .C2(KEYINPUT111), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n554_), .A2(KEYINPUT111), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n760_), .B1(new_n765_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT56), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n550_), .A2(new_n552_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n774_), .A2(KEYINPUT55), .B1(new_n470_), .B2(new_n762_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n774_), .B2(KEYINPUT55), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n777_), .A3(new_n767_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n760_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n771_), .A2(new_n772_), .A3(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n465_), .A2(new_n466_), .A3(new_n560_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n760_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(KEYINPUT112), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n448_), .A2(new_n454_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n449_), .B1(new_n786_), .B2(KEYINPUT113), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n448_), .A2(new_n788_), .A3(new_n454_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n449_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n426_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n785_), .B(new_n463_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n463_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT114), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n563_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n615_), .B1(new_n784_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT57), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n780_), .A2(new_n783_), .B1(new_n563_), .B2(new_n797_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT115), .B(new_n802_), .C1(new_n803_), .C2(new_n615_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n771_), .A2(new_n779_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n561_), .B1(new_n793_), .B2(new_n796_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT116), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n604_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n805_), .A2(new_n806_), .A3(new_n811_), .A4(KEYINPUT58), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n801_), .A2(new_n804_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n759_), .B1(new_n582_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n420_), .A2(new_n384_), .ZN(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n817_));
  OR3_X1    g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n583_), .B1(new_n814_), .B2(KEYINPUT117), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n801_), .A2(new_n820_), .A3(new_n813_), .A4(new_n804_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n759_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT59), .B1(new_n822_), .B2(new_n816_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n818_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n467_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n822_), .A2(new_n816_), .ZN(new_n826_));
  INV_X1    g625(.A(G113gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n701_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(G1340gat));
  INV_X1    g628(.A(G120gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n566_), .B2(KEYINPUT60), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n826_), .B(new_n831_), .C1(KEYINPUT60), .C2(new_n830_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT119), .B1(new_n824_), .B2(new_n566_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G120gat), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n824_), .A2(KEYINPUT119), .A3(new_n566_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n832_), .B1(new_n834_), .B2(new_n835_), .ZN(G1341gat));
  OAI21_X1  g635(.A(G127gat), .B1(new_n824_), .B2(new_n582_), .ZN(new_n837_));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n826_), .A2(new_n838_), .A3(new_n583_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1342gat));
  AOI21_X1  g639(.A(G134gat), .B1(new_n826_), .B2(new_n615_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n824_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT120), .B(G134gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n604_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n842_), .B2(new_n844_), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n814_), .A2(KEYINPUT117), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n582_), .A3(new_n821_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n759_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850_));
  NOR4_X1   g649(.A1(new_n413_), .A2(new_n285_), .A3(new_n421_), .A4(new_n415_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n851_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT121), .B1(new_n822_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n701_), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT122), .B(G141gat), .Z(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1344gat));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n567_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g659(.A1(new_n855_), .A2(new_n583_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  AOI21_X1  g663(.A(G162gat), .B1(new_n855_), .B2(new_n615_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n604_), .A2(new_n203_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n855_), .A2(new_n866_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n615_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n870_), .B(KEYINPUT123), .C1(G162gat), .C2(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n869_), .A2(new_n873_), .ZN(G1347gat));
  NAND2_X1  g673(.A1(new_n421_), .A2(new_n415_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n414_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n657_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n815_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n701_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G169gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT124), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n879_), .A2(new_n882_), .A3(G169gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(KEYINPUT62), .A3(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n878_), .B(KEYINPUT125), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n346_), .A3(new_n701_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n884_), .B(new_n886_), .C1(KEYINPUT62), .C2(new_n881_), .ZN(G1348gat));
  NOR2_X1   g686(.A1(new_n822_), .A2(new_n391_), .ZN(new_n888_));
  AND4_X1   g687(.A1(G176gat), .A2(new_n888_), .A3(new_n567_), .A4(new_n876_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n885_), .A2(new_n567_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n315_), .ZN(G1349gat));
  NOR2_X1   g690(.A1(new_n582_), .A2(new_n328_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n888_), .A2(new_n583_), .A3(new_n876_), .ZN(new_n893_));
  INV_X1    g692(.A(G183gat), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n885_), .A2(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1350gat));
  NAND3_X1  g694(.A1(new_n885_), .A2(new_n341_), .A3(new_n615_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n604_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n885_), .A2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n329_), .ZN(G1351gat));
  NOR4_X1   g698(.A1(new_n822_), .A2(new_n285_), .A3(new_n413_), .A4(new_n875_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n701_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT126), .B(G197gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1352gat));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G204gat), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT127), .B(G204gat), .Z(new_n906_));
  NAND2_X1  g705(.A1(new_n900_), .A2(new_n567_), .ZN(new_n907_));
  MUX2_X1   g706(.A(new_n905_), .B(new_n906_), .S(new_n907_), .Z(G1353gat));
  NAND2_X1  g707(.A1(new_n900_), .A2(new_n583_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  AND2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n909_), .B2(new_n910_), .ZN(G1354gat));
  INV_X1    g712(.A(G218gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n900_), .A2(new_n914_), .A3(new_n615_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n900_), .A2(new_n897_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n914_), .ZN(G1355gat));
endmodule


