//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_;
  INV_X1    g000(.A(G106gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT3), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT2), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n207_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(KEYINPUT1), .B2(new_n208_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(KEYINPUT1), .B2(new_n208_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n203_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(new_n205_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT86), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n211_), .A2(new_n215_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(KEYINPUT29), .A3(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G197gat), .B(G204gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT21), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G211gat), .B(G218gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n223_), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT89), .B1(new_n224_), .B2(new_n225_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT89), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n230_), .B2(new_n227_), .ZN(new_n231_));
  INV_X1    g030(.A(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT88), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(G228gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(G228gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n232_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n221_), .A2(new_n231_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G78gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT29), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n216_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n227_), .A2(new_n230_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n237_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n239_), .A2(new_n240_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n240_), .B1(new_n239_), .B2(new_n245_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n202_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n239_), .A2(new_n245_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G78gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n239_), .A2(new_n240_), .A3(new_n245_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(G106gat), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(new_n252_), .A3(KEYINPUT87), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n217_), .A2(new_n220_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n241_), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT28), .Z(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G22gat), .B(G50gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n256_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n259_), .A2(new_n248_), .A3(new_n252_), .A4(KEYINPUT87), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n257_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n260_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n258_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G1gat), .B(G29gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G85gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT0), .B(G57gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT85), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G113gat), .B(G120gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n217_), .A2(new_n220_), .A3(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT4), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n216_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n274_), .A2(KEYINPUT4), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G225gat), .A2(G233gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n276_), .A2(KEYINPUT93), .A3(new_n279_), .A4(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n274_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n275_), .A2(new_n280_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT93), .B1(new_n285_), .B2(new_n279_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n269_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n279_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT93), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n290_), .A2(new_n268_), .A3(new_n283_), .A4(new_n282_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n293_));
  INV_X1    g092(.A(G169gat), .ZN(new_n294_));
  INV_X1    g093(.A(G176gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT22), .B(G169gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(new_n295_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT23), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n300_), .B(KEYINPUT81), .Z(new_n301_));
  INV_X1    g100(.A(KEYINPUT23), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(G183gat), .A3(G190gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n298_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n296_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT25), .B(G183gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT26), .B(G190gat), .ZN(new_n312_));
  AOI211_X1 g111(.A(new_n308_), .B(new_n310_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n300_), .A2(new_n303_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n307_), .A2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT20), .B1(new_n231_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n313_), .B1(new_n304_), .B2(new_n301_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n306_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n298_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n320_), .B2(new_n298_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n231_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n231_), .A2(KEYINPUT92), .A3(new_n323_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n317_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n293_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n317_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n327_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT92), .B1(new_n231_), .B2(new_n323_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n331_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(KEYINPUT95), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT91), .ZN(new_n339_));
  INV_X1    g138(.A(new_n316_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n244_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n231_), .A2(new_n316_), .A3(KEYINPUT91), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n343_));
  INV_X1    g142(.A(new_n323_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n343_), .B1(new_n344_), .B2(new_n244_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n332_), .B(new_n338_), .C1(new_n337_), .C2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT18), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G64gat), .B(G92gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT32), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n346_), .A2(new_n337_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n333_), .B(new_n331_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT94), .B1(new_n357_), .B2(new_n353_), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n357_), .A2(KEYINPUT94), .A3(new_n353_), .ZN(new_n359_));
  AND4_X1   g158(.A1(new_n292_), .A2(new_n354_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n351_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n355_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n276_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n274_), .A2(new_n278_), .A3(new_n281_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n269_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n284_), .A2(new_n286_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n268_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n291_), .A2(KEYINPUT33), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n367_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n261_), .B(new_n264_), .C1(new_n360_), .C2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n292_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n347_), .A2(new_n361_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n363_), .A2(KEYINPUT27), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n362_), .A2(new_n363_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n375_), .A2(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n257_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n258_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n374_), .B(new_n379_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n373_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT83), .B(G43gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT31), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n323_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G71gat), .B(G99gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT84), .ZN(new_n390_));
  INV_X1    g189(.A(G15gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n388_), .A2(new_n394_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n277_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n277_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n386_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n273_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(new_n396_), .A3(new_n277_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n385_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n380_), .A2(new_n381_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n292_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(KEYINPUT96), .A3(new_n379_), .A4(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n264_), .A2(new_n379_), .A3(new_n261_), .A4(new_n406_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT96), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n383_), .A2(new_n404_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G29gat), .B(G36gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G43gat), .B(G50gat), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G43gat), .B(G50gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT15), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G15gat), .B(G22gat), .ZN(new_n420_));
  INV_X1    g219(.A(G1gat), .ZN(new_n421_));
  INV_X1    g220(.A(G8gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT14), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G1gat), .B(G8gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n419_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n418_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G229gat), .A2(G233gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n426_), .B(new_n428_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G113gat), .B(G141gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G169gat), .B(G197gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n436_), .B(new_n437_), .Z(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n431_), .A2(new_n434_), .A3(new_n438_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(KEYINPUT80), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n443_), .A3(new_n439_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G232gat), .A2(G233gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT35), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n419_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G85gat), .A2(G92gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT7), .ZN(new_n458_));
  INV_X1    g257(.A(G99gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n202_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n462_), .B1(KEYINPUT67), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT67), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n457_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT8), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT66), .ZN(new_n473_));
  INV_X1    g272(.A(G85gat), .ZN(new_n474_));
  INV_X1    g273(.A(G92gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n472_), .A3(new_n453_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n461_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  AOI211_X1 g279(.A(new_n473_), .B(new_n477_), .C1(new_n480_), .C2(new_n467_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n465_), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n460_), .B(new_n461_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n477_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT66), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  OAI22_X1  g285(.A1(new_n471_), .A2(new_n472_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT71), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT10), .B(G99gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n490_), .ZN(new_n492_));
  AOI21_X1  g291(.A(G106gat), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n476_), .A2(KEYINPUT9), .A3(new_n453_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n453_), .A2(KEYINPUT9), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n467_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n488_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n489_), .B(KEYINPUT65), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT71), .B(new_n498_), .C1(new_n499_), .C2(G106gat), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n487_), .A2(KEYINPUT70), .B1(new_n497_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n467_), .A2(KEYINPUT67), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(new_n470_), .A3(new_n480_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n456_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT8), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n464_), .A2(new_n466_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n485_), .B1(new_n506_), .B2(new_n462_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n473_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n484_), .A2(KEYINPUT66), .A3(new_n485_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT70), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n505_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n452_), .B1(new_n501_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n449_), .A2(new_n450_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n487_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(new_n428_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n451_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n481_), .A2(new_n486_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n472_), .B1(new_n503_), .B2(new_n456_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT70), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n497_), .A2(new_n500_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n512_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n419_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n451_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n493_), .A2(new_n496_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n526_), .A2(new_n418_), .B1(new_n450_), .B2(new_n449_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(new_n524_), .A3(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n517_), .A2(KEYINPUT75), .A3(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G190gat), .B(G218gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT36), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n517_), .A2(KEYINPUT75), .A3(new_n528_), .A4(new_n533_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n532_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT36), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n517_), .B2(new_n528_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT37), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n542_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT11), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT68), .B(G71gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G78gat), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n550_), .B(KEYINPUT69), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT11), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n426_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n561_), .B(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT77), .ZN(new_n566_));
  XOR2_X1   g365(.A(G183gat), .B(G211gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(KEYINPUT17), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(KEYINPUT17), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n564_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n573_), .B1(new_n571_), .B2(new_n564_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT78), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n549_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT79), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT64), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n561_), .A2(new_n526_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n561_), .A2(new_n526_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n580_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n556_), .A2(new_n560_), .A3(KEYINPUT12), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n522_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT12), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n561_), .B2(new_n526_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n580_), .B1(new_n561_), .B2(new_n526_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n584_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n591_), .A2(new_n596_), .ZN(new_n599_));
  AND2_X1   g398(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n600_));
  NOR2_X1   g399(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n598_), .B(new_n599_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n591_), .A2(new_n596_), .ZN(new_n603_));
  OAI22_X1  g402(.A1(new_n603_), .A2(new_n597_), .B1(KEYINPUT72), .B2(KEYINPUT13), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT73), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR4_X1   g406(.A1(new_n411_), .A2(new_n446_), .A3(new_n578_), .A4(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n421_), .A3(new_n292_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT38), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n605_), .A2(new_n445_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n383_), .A2(new_n404_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n407_), .A2(new_n410_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n544_), .B(KEYINPUT97), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT98), .B1(new_n411_), .B2(new_n616_), .ZN(new_n619_));
  AOI211_X1 g418(.A(new_n576_), .B(new_n611_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(new_n292_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n610_), .B1(new_n621_), .B2(new_n421_), .ZN(G1324gat));
  INV_X1    g421(.A(new_n379_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n608_), .A2(new_n422_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n623_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n626_), .B2(G8gat), .ZN(new_n627_));
  AOI211_X1 g426(.A(KEYINPUT39), .B(new_n422_), .C1(new_n620_), .C2(new_n623_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n624_), .B(new_n630_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1325gat));
  INV_X1    g433(.A(new_n404_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n608_), .A2(new_n391_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n620_), .A2(new_n635_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT41), .B1(new_n637_), .B2(G15gat), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n639_), .B(new_n391_), .C1(new_n620_), .C2(new_n635_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT100), .B(new_n636_), .C1(new_n638_), .C2(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1326gat));
  INV_X1    g444(.A(G22gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n405_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n620_), .B2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT42), .Z(new_n649_));
  NAND3_X1  g448(.A1(new_n608_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1327gat));
  NOR2_X1   g450(.A1(new_n546_), .A2(new_n547_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT37), .B(new_n542_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT43), .B1(new_n411_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n407_), .A2(new_n410_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n635_), .B1(new_n373_), .B2(new_n382_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n656_), .B(new_n549_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n611_), .A2(new_n575_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(KEYINPUT101), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(KEYINPUT101), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT44), .B1(new_n660_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n667_), .B(new_n664_), .C1(new_n655_), .C2(new_n659_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n666_), .A2(new_n668_), .A3(new_n374_), .ZN(new_n669_));
  INV_X1    g468(.A(G29gat), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n575_), .A2(new_n546_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n605_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n614_), .A2(new_n445_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n292_), .A2(new_n670_), .ZN(new_n674_));
  OAI22_X1  g473(.A1(new_n669_), .A2(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT102), .ZN(G1328gat));
  NAND2_X1  g475(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n666_), .A2(new_n668_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n623_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n379_), .A2(G36gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT103), .B1(new_n673_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n673_), .A2(KEYINPUT103), .A3(new_n686_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n684_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n689_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(KEYINPUT45), .A3(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n677_), .B(new_n680_), .C1(new_n683_), .C2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n666_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n660_), .A2(KEYINPUT44), .A3(new_n665_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n623_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n690_), .A2(new_n692_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n678_), .A4(new_n679_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n694_), .A2(new_n700_), .ZN(G1329gat));
  INV_X1    g500(.A(new_n673_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G43gat), .B1(new_n702_), .B2(new_n635_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n635_), .A2(G43gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n682_), .B2(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g505(.A(G50gat), .B1(new_n702_), .B2(new_n647_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n647_), .A2(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n682_), .B2(new_n708_), .ZN(G1331gat));
  NOR4_X1   g508(.A1(new_n411_), .A2(new_n605_), .A3(new_n578_), .A4(new_n445_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n292_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT105), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n575_), .A2(new_n446_), .ZN(new_n713_));
  AOI211_X1 g512(.A(new_n606_), .B(new_n713_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(G57gat), .A3(new_n292_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1332gat));
  NOR2_X1   g515(.A1(new_n379_), .A2(G64gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT106), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n710_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n714_), .A2(new_n623_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G64gat), .ZN(new_n722_));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT48), .B(new_n723_), .C1(new_n714_), .C2(new_n623_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n719_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT107), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n719_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n710_), .A2(new_n730_), .A3(new_n635_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n714_), .B2(new_n635_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n732_), .A2(new_n733_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1334gat));
  AOI21_X1  g535(.A(new_n240_), .B1(new_n714_), .B2(new_n647_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n710_), .A2(new_n240_), .A3(new_n647_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1335gat));
  NOR3_X1   g540(.A1(new_n605_), .A2(new_n575_), .A3(new_n445_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n655_), .B2(new_n659_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n374_), .ZN(new_n746_));
  AND4_X1   g545(.A1(new_n614_), .A2(new_n446_), .A3(new_n607_), .A4(new_n671_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n474_), .A3(new_n292_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1336gat));
  OAI21_X1  g548(.A(G92gat), .B1(new_n745_), .B2(new_n379_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(new_n475_), .A3(new_n623_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1337gat));
  AOI21_X1  g551(.A(new_n459_), .B1(new_n744_), .B2(new_n635_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n404_), .A2(new_n499_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n747_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n755_), .B(new_n756_), .Z(G1338gat));
  NAND3_X1  g556(.A1(new_n747_), .A2(new_n202_), .A3(new_n647_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n744_), .A2(new_n647_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G106gat), .ZN(new_n761_));
  AOI211_X1 g560(.A(KEYINPUT52), .B(new_n202_), .C1(new_n744_), .C2(new_n647_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g563(.A1(new_n374_), .A2(new_n404_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n405_), .A2(new_n379_), .A3(new_n765_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n654_), .A2(new_n575_), .A3(new_n605_), .A4(new_n446_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n445_), .A2(new_n599_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n586_), .A2(new_n581_), .A3(new_n588_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n580_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n590_), .A2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n586_), .A2(KEYINPUT55), .A3(new_n588_), .A4(new_n589_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n595_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n595_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n770_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n438_), .B1(new_n432_), .B2(new_n430_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n427_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n441_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n546_), .B1(new_n781_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n445_), .A2(new_n599_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n595_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n595_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n790_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n441_), .B(new_n784_), .C1(new_n603_), .C2(new_n597_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(KEYINPUT57), .A3(new_n546_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n789_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n779_), .A2(new_n780_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n603_), .A2(new_n785_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT58), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT112), .B1(new_n800_), .B2(new_n654_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(KEYINPUT58), .A3(new_n799_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n804_), .A2(new_n805_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n797_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT113), .B(new_n769_), .C1(new_n809_), .C2(new_n575_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n805_), .A2(new_n804_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n549_), .A3(new_n807_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n801_), .A2(new_n802_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n795_), .B2(new_n546_), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n788_), .B(new_n544_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n575_), .B1(new_n814_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n768_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n767_), .B(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n811_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n766_), .B1(new_n810_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(G113gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n445_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n818_), .A2(new_n820_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n825_), .A2(KEYINPUT59), .A3(new_n766_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n766_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n814_), .A2(new_n817_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n576_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT113), .B1(new_n829_), .B2(new_n769_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n818_), .A2(new_n820_), .A3(new_n811_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(KEYINPUT59), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT114), .B1(new_n822_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n826_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n837_), .A2(new_n445_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n824_), .B1(new_n838_), .B2(new_n823_), .ZN(G1340gat));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n836_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n826_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n607_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n837_), .A2(KEYINPUT115), .A3(new_n607_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(G120gat), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n605_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n822_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n847_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(G1341gat));
  AOI21_X1  g649(.A(G127gat), .B1(new_n822_), .B2(new_n575_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n575_), .A2(G127gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT116), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n837_), .B2(new_n853_), .ZN(G1342gat));
  INV_X1    g653(.A(G134gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(new_n837_), .B2(new_n549_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n822_), .A2(new_n855_), .A3(new_n616_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT117), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n654_), .B(new_n826_), .C1(new_n834_), .C2(new_n836_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n860_), .B(new_n857_), .C1(new_n861_), .C2(new_n855_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n405_), .A2(new_n635_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n623_), .A2(new_n374_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n864_), .B(new_n865_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n864_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n810_), .B2(new_n821_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT118), .A3(new_n865_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n445_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n872_), .B2(new_n607_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI211_X1 g676(.A(KEYINPUT120), .B(new_n606_), .C1(new_n868_), .C2(new_n871_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT119), .B(G148gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n877_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n880_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1345gat));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n872_), .B2(new_n575_), .ZN(new_n886_));
  AOI211_X1 g685(.A(KEYINPUT121), .B(new_n576_), .C1(new_n868_), .C2(new_n871_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n886_), .A2(new_n887_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n810_), .A2(new_n821_), .ZN(new_n891_));
  AND4_X1   g690(.A1(KEYINPUT118), .A2(new_n891_), .A3(new_n864_), .A4(new_n865_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT118), .B1(new_n870_), .B2(new_n865_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n575_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT121), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n872_), .A2(new_n885_), .A3(new_n575_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n888_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n890_), .A2(new_n897_), .ZN(G1346gat));
  INV_X1    g697(.A(G162gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n872_), .A2(new_n899_), .A3(new_n616_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n654_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1347gat));
  INV_X1    g701(.A(new_n825_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n379_), .A2(new_n292_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n635_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n446_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n906_), .A2(KEYINPUT122), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(KEYINPUT122), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n647_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n294_), .B1(new_n903_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(KEYINPUT62), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n825_), .A2(new_n647_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(new_n297_), .A3(new_n906_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n915_));
  OAI211_X1 g714(.A(new_n912_), .B(new_n914_), .C1(new_n910_), .C2(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT124), .ZN(G1348gat));
  NAND3_X1  g716(.A1(new_n913_), .A2(new_n635_), .A3(new_n904_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n295_), .B1(new_n918_), .B2(new_n605_), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT125), .Z(new_n920_));
  AOI21_X1  g719(.A(new_n647_), .B1(new_n810_), .B2(new_n821_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n606_), .A2(new_n905_), .A3(new_n295_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(G1349gat));
  INV_X1    g722(.A(new_n311_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n905_), .A2(new_n576_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n913_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT126), .ZN(new_n927_));
  AOI21_X1  g726(.A(G183gat), .B1(new_n921_), .B2(new_n925_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(KEYINPUT127), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n918_), .B2(new_n654_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n616_), .A2(new_n312_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n918_), .B2(new_n932_), .ZN(G1351gat));
  AND2_X1   g732(.A1(new_n870_), .A2(new_n904_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n445_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n607_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g737(.A(new_n576_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n934_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  XOR2_X1   g740(.A(new_n940_), .B(new_n941_), .Z(G1354gat));
  INV_X1    g741(.A(G218gat), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n934_), .A2(new_n943_), .A3(new_n616_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n934_), .A2(new_n549_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n943_), .ZN(G1355gat));
endmodule


