//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(G15gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G71gat), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT82), .B(G43gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G169gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT79), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT22), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT79), .B1(new_n211_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n209_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(G176gat), .B1(new_n211_), .B2(KEYINPUT79), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT22), .B(G169gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n219_), .B(KEYINPUT80), .C1(KEYINPUT79), .C2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G183gat), .A3(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n226_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n218_), .A2(new_n221_), .A3(new_n223_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT78), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n225_), .A2(new_n227_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(KEYINPUT24), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n235_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n225_), .A2(new_n227_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n241_), .B(KEYINPUT78), .C1(KEYINPUT24), .C2(new_n238_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT25), .B(G183gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT26), .B(G190gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n222_), .A2(new_n237_), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n243_), .A2(new_n244_), .B1(new_n245_), .B2(KEYINPUT24), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n240_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n234_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT30), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT83), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n208_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n249_), .B(KEYINPUT83), .Z(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n252_), .B2(new_n208_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G127gat), .B(G134gat), .Z(new_n254_));
  XOR2_X1   g053(.A(G113gat), .B(G120gat), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G127gat), .B(G134gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n256_), .A2(KEYINPUT84), .A3(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n253_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n253_), .A2(new_n267_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G85gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT0), .B(G57gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  NAND2_X1  g073(.A1(G225gat), .A2(G233gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT2), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(G141gat), .A3(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT3), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n281_), .A2(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT87), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT87), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n289_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT88), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n286_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n279_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n276_), .A2(KEYINPUT1), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n276_), .B1(new_n278_), .B2(KEYINPUT1), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT86), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(KEYINPUT86), .B(new_n276_), .C1(new_n278_), .C2(KEYINPUT1), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n280_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(new_n285_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n295_), .A2(new_n304_), .B1(new_n263_), .B2(new_n262_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n275_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n279_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n288_), .A2(new_n290_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n285_), .A2(new_n284_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n282_), .B1(G141gat), .B2(G148gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n280_), .A2(KEYINPUT2), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT88), .B1(new_n309_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n286_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n308_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n301_), .A2(new_n303_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n264_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n295_), .A2(new_n260_), .A3(new_n304_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT4), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n307_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n319_), .A3(new_n275_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n274_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n318_), .A2(KEYINPUT4), .A3(new_n319_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n275_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n318_), .B2(KEYINPUT4), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n322_), .B(new_n274_), .C1(new_n325_), .C2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n270_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n332_));
  NAND2_X1  g131(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n334_), .A2(new_n335_), .A3(G197gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT21), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(G197gat), .B2(G204gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n332_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G197gat), .ZN(new_n341_));
  OR2_X1    g140(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n333_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n337_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n333_), .ZN(new_n347_));
  OAI211_X1 g146(.A(KEYINPUT90), .B(new_n338_), .C1(new_n347_), .C2(G197gat), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n340_), .A2(new_n345_), .A3(new_n346_), .A4(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n343_), .A2(new_n344_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT91), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n337_), .B1(new_n346_), .B2(new_n351_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n350_), .B(new_n352_), .C1(new_n351_), .C2(new_n346_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n211_), .A2(new_n216_), .A3(new_n213_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n223_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n231_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n245_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n243_), .A2(new_n244_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n237_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n229_), .A2(new_n230_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n358_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n354_), .A2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n234_), .A2(new_n349_), .A3(new_n247_), .A4(new_n353_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(KEYINPUT20), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT19), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n248_), .A2(new_n354_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n248_), .B2(new_n354_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n356_), .A2(new_n357_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n365_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n380_), .A2(KEYINPUT95), .A3(new_n353_), .A4(new_n349_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n354_), .B2(new_n366_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n371_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n372_), .B1(new_n376_), .B2(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(G8gat), .B(G36gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n387_), .A2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n372_), .B(new_n392_), .C1(new_n376_), .C2(new_n386_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT27), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT101), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(KEYINPUT101), .A3(new_n397_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT20), .B1(new_n354_), .B2(new_n366_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n371_), .B1(new_n376_), .B2(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n369_), .A2(new_n371_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n393_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n395_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(new_n397_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n400_), .A2(new_n401_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n295_), .A2(new_n304_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT29), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n354_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(G228gat), .A3(G233gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n416_), .A3(new_n354_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n411_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n415_), .A2(new_n417_), .A3(new_n411_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n412_), .A2(KEYINPUT29), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G22gat), .B(G50gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT28), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n422_), .B(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n418_), .B2(KEYINPUT92), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n419_), .A2(KEYINPUT92), .A3(new_n420_), .A4(new_n425_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n409_), .A2(KEYINPUT102), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT102), .ZN(new_n431_));
  INV_X1    g230(.A(new_n429_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n408_), .A2(new_n406_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT101), .B1(new_n396_), .B2(new_n397_), .ZN(new_n434_));
  AOI211_X1 g233(.A(new_n399_), .B(KEYINPUT27), .C1(new_n394_), .C2(new_n395_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n431_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n331_), .B1(new_n430_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n381_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n248_), .A2(new_n354_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT94), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n248_), .A2(new_n354_), .A3(new_n373_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n392_), .B1(new_n445_), .B2(new_n372_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n439_), .B1(new_n446_), .B2(new_n407_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n318_), .A2(new_n319_), .A3(new_n326_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n274_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n326_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n320_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT98), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(KEYINPUT33), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n328_), .A2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n321_), .A2(new_n322_), .A3(new_n274_), .A4(new_n454_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n452_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n394_), .A2(KEYINPUT97), .A3(new_n395_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n447_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n392_), .A2(KEYINPUT32), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n445_), .A2(new_n461_), .A3(new_n372_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n321_), .A2(new_n322_), .A3(new_n274_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n323_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT99), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n461_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n405_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT99), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n329_), .A2(new_n468_), .A3(new_n469_), .A4(new_n462_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n460_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n429_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT100), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n429_), .A2(new_n329_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n472_), .A2(new_n473_), .B1(new_n409_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n471_), .A2(KEYINPUT100), .A3(new_n429_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n270_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n438_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G85gat), .A2(G92gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT69), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT8), .B1(new_n483_), .B2(KEYINPUT68), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT67), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n491_));
  OAI22_X1  g290(.A1(new_n490_), .A2(new_n491_), .B1(G99gat), .B2(G106gat), .ZN(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n205_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n494_), .B2(new_n490_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n483_), .B1(new_n487_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n484_), .A2(new_n496_), .ZN(new_n497_));
  OAI221_X1 g296(.A(new_n483_), .B1(KEYINPUT68), .B2(KEYINPUT8), .C1(new_n487_), .C2(new_n495_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n486_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n485_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n485_), .A2(new_n499_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  AOI22_X1  g301(.A1(new_n500_), .A2(new_n501_), .B1(new_n493_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT64), .B(G85gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT9), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(G92gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n480_), .A2(KEYINPUT9), .A3(new_n481_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n503_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n497_), .A2(new_n498_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n517_));
  XOR2_X1   g316(.A(G71gat), .B(G78gat), .Z(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n517_), .A2(new_n518_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT70), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n513_), .A2(new_n520_), .A3(new_n519_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n525_), .B(new_n527_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT71), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n503_), .B(new_n529_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n506_), .A2(new_n508_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT65), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n509_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n529_), .B1(new_n534_), .B2(new_n503_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n498_), .B(new_n497_), .C1(new_n531_), .C2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT12), .B1(new_n521_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n538_), .B1(new_n537_), .B2(new_n521_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n536_), .A2(new_n539_), .B1(new_n514_), .B2(new_n521_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n524_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n526_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n528_), .A2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G120gat), .B(G148gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n528_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n553_), .A2(KEYINPUT13), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(KEYINPUT13), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G29gat), .B(G36gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT75), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561_));
  INV_X1    g360(.A(G1gat), .ZN(new_n562_));
  INV_X1    g361(.A(G8gat), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT14), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G1gat), .B(G8gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n560_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n560_), .B(KEYINPUT15), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n567_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n569_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n567_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n560_), .B2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n570_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G169gat), .B(G197gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(KEYINPUT77), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n576_), .B(new_n580_), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n556_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n479_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT34), .Z(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n536_), .A2(new_n571_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n514_), .A2(new_n560_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n589_), .A2(new_n590_), .A3(new_n588_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n595_), .B(KEYINPUT36), .Z(new_n599_));
  INV_X1    g398(.A(new_n597_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n599_), .B1(new_n600_), .B2(new_n591_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n601_), .A3(KEYINPUT76), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT37), .Z(new_n603_));
  XNOR2_X1  g402(.A(new_n521_), .B(new_n567_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(G127gat), .B(G155gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT16), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT17), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n537_), .A2(KEYINPUT17), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n612_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n606_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n610_), .A2(new_n613_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n606_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n603_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n583_), .A2(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n620_), .A2(G1gat), .A3(new_n330_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT38), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT38), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n598_), .A2(new_n601_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n479_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n582_), .A2(new_n618_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n330_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n622_), .A2(new_n623_), .A3(new_n631_), .ZN(G1324gat));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n436_), .A3(new_n629_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n563_), .B1(KEYINPUT104), .B2(KEYINPUT39), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n436_), .A2(new_n563_), .ZN(new_n638_));
  OAI22_X1  g437(.A1(new_n636_), .A2(new_n637_), .B1(new_n620_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n639_), .B(new_n640_), .Z(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n630_), .B2(new_n478_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT41), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n620_), .A2(G15gat), .A3(new_n478_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1326gat));
  OAI21_X1  g444(.A(G22gat), .B1(new_n630_), .B2(new_n429_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT42), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n429_), .A2(G22gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n620_), .B2(new_n648_), .ZN(G1327gat));
  INV_X1    g448(.A(new_n627_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n618_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n583_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G29gat), .B1(new_n654_), .B2(new_n329_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n270_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n656_), .B(new_n603_), .C1(new_n657_), .C2(new_n438_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT106), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n430_), .A2(new_n437_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n331_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n476_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n436_), .A2(new_n429_), .A3(new_n329_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT100), .B1(new_n471_), .B2(new_n429_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n666_), .B2(new_n270_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n656_), .A4(new_n603_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n602_), .B(KEYINPUT37), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT43), .B1(new_n479_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n659_), .A2(new_n669_), .A3(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n582_), .A2(new_n651_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT44), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n673_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n672_), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n673_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n329_), .A2(G29gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n655_), .B1(new_n679_), .B2(new_n680_), .ZN(G1328gat));
  INV_X1    g480(.A(G36gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n436_), .A2(new_n682_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n653_), .A2(KEYINPUT108), .A3(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT108), .B1(new_n653_), .B2(new_n683_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(KEYINPUT45), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT45), .B1(new_n684_), .B2(new_n685_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI211_X1 g488(.A(new_n409_), .B(new_n674_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n689_), .B(KEYINPUT46), .C1(new_n690_), .C2(new_n682_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n677_), .A2(new_n678_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n674_), .A2(new_n409_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n682_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n684_), .A2(new_n685_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n686_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n692_), .B1(new_n695_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n691_), .A2(new_n700_), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n270_), .A2(G43gat), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n674_), .B(new_n702_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G43gat), .B1(new_n654_), .B2(new_n270_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT47), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n679_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708_));
  INV_X1    g507(.A(new_n704_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n705_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n654_), .B2(new_n432_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n432_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n679_), .B2(new_n713_), .ZN(G1331gat));
  NOR3_X1   g513(.A1(new_n479_), .A2(new_n581_), .A3(new_n556_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n619_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n330_), .B1(new_n716_), .B2(KEYINPUT109), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(KEYINPUT109), .B2(new_n716_), .ZN(new_n718_));
  INV_X1    g517(.A(G57gat), .ZN(new_n719_));
  INV_X1    g518(.A(new_n556_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n581_), .A2(new_n618_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n628_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n330_), .A2(new_n719_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n718_), .A2(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n722_), .B2(new_n436_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT48), .Z(new_n727_));
  NAND2_X1  g526(.A1(new_n436_), .A2(new_n725_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n716_), .B2(new_n728_), .ZN(G1333gat));
  OR3_X1    g528(.A1(new_n716_), .A2(G71gat), .A3(new_n478_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n722_), .A2(new_n270_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT49), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(G71gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n731_), .B2(G71gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT110), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n722_), .B2(new_n432_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT50), .Z(new_n739_));
  NOR2_X1   g538(.A1(new_n429_), .A2(G78gat), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT111), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n716_), .B2(new_n741_), .ZN(G1335gat));
  NAND2_X1  g541(.A1(new_n715_), .A2(new_n652_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n715_), .A2(KEYINPUT112), .A3(new_n652_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n329_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n556_), .A2(new_n651_), .A3(new_n581_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n672_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n329_), .A2(new_n504_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT113), .Z(new_n752_));
  AOI21_X1  g551(.A(new_n748_), .B1(new_n750_), .B2(new_n752_), .ZN(G1336gat));
  INV_X1    g552(.A(G92gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n747_), .A2(new_n754_), .A3(new_n436_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n750_), .A2(new_n436_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n754_), .ZN(G1337gat));
  NAND2_X1  g556(.A1(new_n270_), .A2(new_n502_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT114), .B1(new_n747_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  AOI211_X1 g560(.A(new_n761_), .B(new_n758_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n750_), .A2(new_n270_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(new_n205_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT51), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767_));
  OAI221_X1 g566(.A(new_n767_), .B1(new_n764_), .B2(new_n205_), .C1(new_n760_), .C2(new_n762_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1338gat));
  NAND3_X1  g568(.A1(new_n747_), .A2(new_n493_), .A3(new_n432_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n672_), .A2(new_n432_), .A3(new_n749_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  AND4_X1   g571(.A1(KEYINPUT115), .A2(new_n771_), .A3(new_n772_), .A4(G106gat), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n493_), .B1(new_n774_), .B2(KEYINPUT52), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n771_), .A2(new_n775_), .B1(KEYINPUT115), .B2(new_n772_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n770_), .B1(new_n773_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n770_), .C1(new_n773_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  NAND3_X1  g580(.A1(new_n660_), .A2(new_n270_), .A3(new_n329_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT121), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n526_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n543_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n540_), .A2(KEYINPUT55), .A3(new_n526_), .A4(new_n542_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n549_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n552_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n579_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n576_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n569_), .B1(new_n560_), .B2(new_n574_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n572_), .A2(new_n794_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n568_), .A2(new_n573_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n579_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n793_), .A2(new_n797_), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT56), .B(new_n549_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n791_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n603_), .B(new_n784_), .C1(new_n800_), .C2(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n787_), .A2(new_n788_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n550_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT56), .ZN(new_n806_));
  INV_X1    g605(.A(new_n798_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n789_), .A2(new_n790_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n806_), .A2(new_n552_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n784_), .B1(new_n811_), .B2(new_n603_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n803_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n806_), .A2(new_n581_), .A3(new_n552_), .A4(new_n808_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n553_), .A2(new_n807_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n627_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n816_), .B(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n618_), .B1(new_n813_), .B2(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n721_), .B(KEYINPUT116), .Z(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(new_n670_), .A3(new_n556_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n821_), .A2(new_n670_), .A3(new_n556_), .A4(new_n823_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n820_), .A2(KEYINPUT120), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n603_), .B1(new_n800_), .B2(KEYINPUT58), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT119), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n802_), .A3(new_n801_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n814_), .A2(new_n815_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n818_), .B1(new_n834_), .B2(new_n650_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n627_), .B(new_n817_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n651_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n838_), .B2(new_n827_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n783_), .B1(new_n829_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(G113gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n581_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n820_), .A2(new_n828_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n783_), .B2(KEYINPUT123), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n843_), .B(new_n845_), .C1(KEYINPUT123), .C2(new_n783_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n581_), .B(new_n846_), .C1(new_n840_), .C2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n842_), .B1(new_n849_), .B2(new_n841_), .ZN(G1340gat));
  OAI21_X1  g649(.A(new_n846_), .B1(new_n840_), .B2(new_n847_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G120gat), .B1(new_n851_), .B2(new_n556_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n840_), .ZN(new_n853_));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n556_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(KEYINPUT60), .B2(new_n854_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n852_), .B1(new_n853_), .B2(new_n856_), .ZN(G1341gat));
  INV_X1    g656(.A(G127gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n651_), .B2(KEYINPUT124), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(KEYINPUT124), .B2(new_n858_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n846_), .B(new_n860_), .C1(new_n840_), .C2(new_n847_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n783_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT120), .B1(new_n820_), .B2(new_n828_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n838_), .A2(new_n830_), .A3(new_n827_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n651_), .B(new_n862_), .C1(new_n863_), .C2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n858_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n861_), .A2(KEYINPUT125), .A3(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1342gat));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n840_), .A2(new_n872_), .A3(new_n627_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n603_), .B(new_n846_), .C1(new_n840_), .C2(new_n847_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n875_), .B2(new_n872_), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n270_), .A2(new_n429_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n329_), .A3(new_n409_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n829_), .B2(new_n839_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n581_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n720_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n879_), .A2(new_n886_), .A3(new_n651_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n879_), .B2(new_n651_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n889_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n887_), .A3(new_n884_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1346gat));
  INV_X1    g692(.A(G162gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n879_), .A2(new_n894_), .A3(new_n627_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n879_), .A2(new_n603_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n894_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n331_), .A2(new_n409_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n432_), .B(new_n900_), .C1(new_n820_), .C2(new_n828_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n581_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n898_), .B1(new_n903_), .B2(new_n215_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n220_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n902_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(G1348gat));
  AOI21_X1  g706(.A(G176gat), .B1(new_n901_), .B2(new_n720_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n432_), .B1(new_n829_), .B2(new_n839_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n900_), .A2(new_n213_), .A3(new_n556_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1349gat));
  NAND3_X1  g710(.A1(new_n909_), .A2(new_n651_), .A3(new_n899_), .ZN(new_n912_));
  INV_X1    g711(.A(G183gat), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n618_), .A2(new_n243_), .ZN(new_n914_));
  AOI22_X1  g713(.A1(new_n912_), .A2(new_n913_), .B1(new_n901_), .B2(new_n914_), .ZN(G1350gat));
  NAND2_X1  g714(.A1(new_n901_), .A2(new_n603_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G190gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n901_), .A2(new_n244_), .A3(new_n627_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1351gat));
  NAND3_X1  g718(.A1(new_n877_), .A2(new_n330_), .A3(new_n436_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(new_n829_), .B2(new_n839_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n581_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g722(.A1(new_n921_), .A2(new_n720_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(G204gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n347_), .B2(new_n924_), .ZN(G1353gat));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n927_));
  INV_X1    g726(.A(G211gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n651_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(KEYINPUT127), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n921_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n927_), .A2(new_n928_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1354gat));
  INV_X1    g732(.A(G218gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n921_), .A2(new_n934_), .A3(new_n627_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n921_), .A2(new_n603_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n934_), .ZN(G1355gat));
endmodule


