//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT64), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT7), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G85gat), .B(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n212_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n205_), .B(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n208_), .A2(new_n210_), .A3(new_n219_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n214_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n216_), .B1(new_n223_), .B2(new_n213_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT10), .B(G99gat), .Z(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT65), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229_));
  MUX2_X1   g028(.A(new_n229_), .B(new_n214_), .S(KEYINPUT9), .Z(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n211_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n235_));
  XOR2_X1   g034(.A(G71gat), .B(G78gat), .Z(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n235_), .A2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n224_), .A2(new_n231_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n239_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n241_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n243_), .A2(KEYINPUT67), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n204_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT68), .B(new_n216_), .C1(new_n223_), .C2(new_n213_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n211_), .A2(KEYINPUT66), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n206_), .A3(new_n222_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n213_), .B1(new_n252_), .B2(new_n215_), .ZN(new_n253_));
  AOI211_X1 g052(.A(KEYINPUT8), .B(new_n214_), .C1(new_n206_), .C2(new_n211_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n250_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n231_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n240_), .A2(KEYINPUT12), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n241_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n243_), .A3(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n263_), .A2(new_n204_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G120gat), .B(G148gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n248_), .A2(new_n264_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n270_), .B1(new_n248_), .B2(new_n264_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n275_), .A2(KEYINPUT13), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n275_), .A2(KEYINPUT13), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n274_), .B1(new_n278_), .B2(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G218gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G211gat), .ZN(new_n283_));
  INV_X1    g082(.A(G211gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G218gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT90), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G211gat), .B(G218gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT90), .ZN(new_n290_));
  INV_X1    g089(.A(G197gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT87), .B1(new_n291_), .B2(G204gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT87), .ZN(new_n293_));
  INV_X1    g092(.A(G204gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(G197gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(G204gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n288_), .A2(new_n290_), .A3(KEYINPUT21), .A4(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n299_));
  NAND4_X1  g098(.A1(new_n299_), .A2(new_n292_), .A3(new_n295_), .A4(new_n296_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(G197gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n296_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n286_), .B1(KEYINPUT21), .B2(new_n302_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n300_), .A2(new_n303_), .A3(KEYINPUT89), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT89), .B1(new_n300_), .B2(new_n303_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n298_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307_));
  INV_X1    g106(.A(G141gat), .ZN(new_n308_));
  INV_X1    g107(.A(G148gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT2), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n310_), .A2(new_n313_), .A3(new_n314_), .A4(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n308_), .A2(new_n309_), .A3(KEYINPUT82), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(G141gat), .B2(G148gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n317_), .A2(new_n325_), .A3(new_n318_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n327_), .A2(new_n311_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n320_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT83), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n320_), .A2(new_n329_), .A3(KEYINPUT83), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT29), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n335_), .B(KEYINPUT86), .Z(new_n336_));
  NAND3_X1  g135(.A1(new_n306_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n330_), .A2(KEYINPUT29), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n306_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT91), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AOI211_X1 g140(.A(KEYINPUT91), .B(new_n336_), .C1(new_n306_), .C2(new_n338_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n337_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(KEYINPUT92), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n337_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n298_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n302_), .A2(KEYINPUT21), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n350_), .B(new_n289_), .C1(new_n297_), .C2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n300_), .A2(new_n303_), .A3(KEYINPUT89), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n349_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n338_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT91), .B1(new_n358_), .B2(new_n336_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n339_), .A2(new_n340_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n348_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n345_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n347_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT85), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n332_), .A2(new_n333_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n320_), .A2(KEYINPUT83), .A3(new_n329_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT83), .B1(new_n320_), .B2(new_n329_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n365_), .B(new_n367_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT84), .B1(new_n368_), .B2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G22gat), .B(G50gat), .Z(new_n374_));
  OAI21_X1  g173(.A(new_n367_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT28), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT84), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n371_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n373_), .A2(new_n374_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n374_), .B1(new_n373_), .B2(new_n378_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n364_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n373_), .A2(new_n378_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n374_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(KEYINPUT85), .A3(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n363_), .A2(new_n382_), .A3(new_n386_), .ZN(new_n387_));
  OR3_X1    g186(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n388_));
  AND2_X1   g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT26), .B(G190gat), .ZN(new_n392_));
  INV_X1    g191(.A(G183gat), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n393_), .A2(KEYINPUT25), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(KEYINPUT25), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT78), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n391_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G183gat), .A2(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT79), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(G183gat), .A3(G190gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT23), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT23), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(G183gat), .B2(G190gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n398_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n400_), .A2(new_n402_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT23), .ZN(new_n410_));
  OR2_X1    g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n399_), .A2(new_n404_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G169gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n408_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G227gat), .A2(G233gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n418_), .B(KEYINPUT80), .Z(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT30), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n417_), .B(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G71gat), .B(G99gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G127gat), .B(G134gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G113gat), .B(G120gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT31), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n428_), .B2(new_n427_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G15gat), .B(G43gat), .Z(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n423_), .B(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n385_), .A2(new_n379_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n344_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT93), .B1(new_n361_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT93), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n343_), .A2(new_n437_), .A3(new_n344_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .A4(new_n362_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n387_), .A2(new_n433_), .A3(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G8gat), .B(G36gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT18), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G64gat), .B(G92gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n398_), .A2(new_n407_), .B1(new_n415_), .B2(new_n413_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n356_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n415_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT96), .ZN(new_n450_));
  INV_X1    g249(.A(new_n411_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n406_), .B2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT96), .B(new_n411_), .C1(new_n403_), .C2(new_n405_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n410_), .A2(new_n412_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n391_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n392_), .A2(new_n396_), .A3(new_n394_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n306_), .B1(new_n454_), .B2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n461_));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT95), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n448_), .A2(new_n460_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n452_), .A2(new_n453_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n415_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(new_n356_), .A3(new_n458_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n446_), .B1(new_n306_), .B2(new_n417_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n463_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n445_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n464_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n356_), .B1(new_n467_), .B2(new_n458_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT20), .B1(new_n306_), .B2(new_n417_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n468_), .A2(new_n469_), .A3(new_n463_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n444_), .A3(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n471_), .A2(KEYINPUT27), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT97), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n475_), .A2(KEYINPUT97), .A3(new_n444_), .A4(new_n476_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n475_), .A2(new_n476_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n445_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n479_), .B1(new_n485_), .B2(KEYINPUT27), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G225gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n427_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT98), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n332_), .A2(new_n488_), .A3(new_n489_), .A4(new_n333_), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n369_), .A2(new_n370_), .A3(new_n427_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT98), .B1(new_n488_), .B2(new_n330_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n487_), .B(new_n490_), .C1(new_n491_), .C2(new_n492_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n366_), .A2(KEYINPUT4), .A3(new_n427_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(new_n495_), .B2(KEYINPUT4), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n493_), .B1(new_n496_), .B2(new_n487_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G1gat), .B(G29gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G85gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT0), .B(G57gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n493_), .B(new_n501_), .C1(new_n496_), .C2(new_n487_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n440_), .A2(new_n486_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n387_), .A2(new_n439_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT27), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n478_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n505_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n444_), .A2(KEYINPUT32), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(new_n513_), .B2(new_n483_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n504_), .B2(new_n503_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n503_), .A2(KEYINPUT33), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT33), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n497_), .A2(new_n518_), .A3(new_n502_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n496_), .A2(new_n487_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT99), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n495_), .A2(G225gat), .A3(G233gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n501_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n520_), .B2(KEYINPUT99), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n517_), .A2(new_n519_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n516_), .B1(new_n525_), .B2(new_n485_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n512_), .B1(new_n526_), .B2(new_n507_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n433_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n506_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT76), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G29gat), .B(G36gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT71), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G43gat), .B(G50gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537_));
  INV_X1    g336(.A(G1gat), .ZN(new_n538_));
  INV_X1    g337(.A(G8gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G1gat), .B(G8gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  NOR2_X1   g342(.A1(new_n536_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n535_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n534_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n543_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n532_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n548_), .A2(new_n544_), .A3(new_n532_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n531_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n536_), .A2(KEYINPUT15), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n547_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n548_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n552_), .B1(new_n531_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n552_), .B(new_n563_), .C1(new_n531_), .C2(new_n559_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT77), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n560_), .A2(KEYINPUT77), .A3(new_n564_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n281_), .A2(new_n529_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n257_), .A2(new_n556_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n224_), .A2(new_n231_), .A3(new_n536_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT34), .Z(new_n575_));
  INV_X1    g374(.A(KEYINPUT35), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT72), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT73), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n575_), .A2(new_n576_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n572_), .A2(new_n580_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n581_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT73), .B1(new_n575_), .B2(new_n576_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n256_), .A2(new_n231_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n584_), .B(new_n585_), .C1(new_n586_), .C2(new_n579_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n583_), .A2(new_n587_), .A3(new_n594_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n593_), .A2(new_n595_), .B1(KEYINPUT36), .B2(new_n591_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n593_), .B2(KEYINPUT74), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n600_));
  INV_X1    g399(.A(new_n595_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n594_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n600_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT37), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n599_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n543_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(new_n239_), .ZN(new_n611_));
  XOR2_X1   g410(.A(G127gat), .B(G155gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT16), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT75), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n615_), .A2(new_n616_), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n611_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n608_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n571_), .A2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(KEYINPUT100), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(KEYINPUT100), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n625_), .A2(new_n538_), .A3(new_n505_), .A4(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n622_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n596_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n571_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n538_), .B1(new_n633_), .B2(new_n505_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n629_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n628_), .B2(new_n627_), .ZN(G1324gat));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n486_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(G8gat), .ZN(new_n639_));
  AOI211_X1 g438(.A(KEYINPUT39), .B(new_n539_), .C1(new_n633_), .C2(new_n486_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n625_), .A2(new_n539_), .A3(new_n486_), .A4(new_n626_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(G1325gat));
  INV_X1    g444(.A(G15gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n633_), .B2(new_n433_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT41), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n433_), .A2(new_n646_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n624_), .B2(new_n649_), .ZN(G1326gat));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n633_), .B2(new_n507_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n507_), .A2(new_n651_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT103), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n654_), .B1(new_n624_), .B2(new_n656_), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n630_), .A2(new_n596_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n571_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(G29gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n505_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n607_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n599_), .A2(new_n606_), .A3(KEYINPUT104), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n529_), .B2(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n607_), .A2(KEYINPUT43), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT105), .B1(new_n529_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n607_), .A2(KEYINPUT43), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n521_), .A2(new_n524_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n519_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n518_), .B1(new_n497_), .B2(new_n502_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  OAI22_X1  g474(.A1(new_n675_), .A2(new_n508_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n507_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n433_), .B1(new_n678_), .B2(new_n512_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n670_), .B(new_n671_), .C1(new_n679_), .C2(new_n506_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n667_), .A2(new_n669_), .A3(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n281_), .A2(new_n570_), .A3(new_n630_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT44), .B1(new_n681_), .B2(new_n682_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n511_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n662_), .B1(new_n685_), .B2(new_n661_), .ZN(G1328gat));
  NOR3_X1   g485(.A1(new_n659_), .A2(G36gat), .A3(new_n510_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n683_), .A2(new_n684_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT106), .B1(new_n690_), .B2(new_n486_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n681_), .A2(new_n682_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n682_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n694_), .A2(KEYINPUT106), .A3(new_n486_), .A4(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n689_), .B1(new_n691_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n694_), .A2(new_n486_), .A3(new_n695_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(G36gat), .A3(new_n696_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n707_), .A2(new_n699_), .A3(new_n700_), .A4(new_n689_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n703_), .A2(new_n708_), .ZN(G1329gat));
  NAND3_X1  g508(.A1(new_n690_), .A2(G43gat), .A3(new_n433_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n659_), .A2(new_n528_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(G43gat), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g512(.A(G50gat), .B1(new_n660_), .B2(new_n507_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n507_), .A2(G50gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n690_), .B2(new_n715_), .ZN(G1331gat));
  INV_X1    g515(.A(new_n570_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n529_), .A2(new_n280_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n623_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT108), .Z(new_n720_));
  INV_X1    g519(.A(G57gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n505_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n718_), .A2(new_n632_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n511_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1332gat));
  INV_X1    g525(.A(G64gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n723_), .B2(new_n486_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT109), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n720_), .A2(new_n727_), .A3(new_n486_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(G1333gat));
  INV_X1    g532(.A(G71gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n723_), .B2(new_n433_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT49), .Z(new_n736_));
  NAND2_X1  g535(.A1(new_n433_), .A2(new_n734_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT110), .Z(new_n738_));
  NAND2_X1  g537(.A1(new_n720_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n723_), .B2(new_n507_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT50), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n720_), .A2(new_n741_), .A3(new_n507_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1335gat));
  AND2_X1   g544(.A1(new_n718_), .A2(new_n658_), .ZN(new_n746_));
  INV_X1    g545(.A(G85gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n505_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n280_), .A2(new_n717_), .A3(new_n630_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n681_), .A2(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n511_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n753_), .B2(new_n747_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT112), .ZN(G1336gat));
  INV_X1    g554(.A(G92gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n746_), .A2(new_n756_), .A3(new_n486_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n751_), .A2(new_n752_), .A3(new_n510_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(new_n756_), .ZN(G1337gat));
  NAND2_X1  g558(.A1(new_n750_), .A2(new_n433_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n433_), .A2(new_n225_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n760_), .A2(G99gat), .B1(new_n746_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n681_), .A2(new_n507_), .A3(new_n749_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT115), .B1(new_n765_), .B2(G106gat), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n768_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n746_), .A2(new_n226_), .A3(new_n507_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT114), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n769_), .A2(new_n775_), .A3(new_n770_), .A4(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  AOI21_X1  g576(.A(new_n244_), .B1(new_n261_), .B2(new_n241_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n778_), .A2(KEYINPUT55), .A3(new_n203_), .A4(new_n260_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n263_), .B2(new_n204_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n263_), .A2(new_n204_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n269_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n269_), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n272_), .B(new_n570_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n548_), .A2(new_n544_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT76), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n531_), .B1(new_n790_), .B2(new_n549_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT116), .B1(new_n791_), .B2(new_n563_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n530_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n564_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n559_), .A2(KEYINPUT117), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n557_), .A2(new_n797_), .A3(new_n558_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n531_), .A3(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n792_), .A2(new_n795_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n792_), .A2(new_n795_), .A3(new_n799_), .A4(KEYINPUT118), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n566_), .A3(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(new_n274_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n596_), .B1(new_n788_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n787_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n783_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n269_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n786_), .A3(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n804_), .A2(new_n272_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n607_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n813_), .A3(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT120), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n812_), .A2(new_n813_), .A3(new_n819_), .A4(KEYINPUT58), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n806_), .A2(new_n807_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n808_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(new_n822_), .A3(KEYINPUT121), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n630_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n623_), .A2(new_n280_), .A3(new_n570_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT54), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n440_), .A2(new_n486_), .A3(new_n511_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n622_), .B1(new_n823_), .B2(new_n808_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n829_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n836_), .A2(new_n832_), .ZN(new_n837_));
  OAI22_X1  g636(.A1(new_n831_), .A2(new_n834_), .B1(new_n837_), .B2(new_n833_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n570_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n837_), .ZN(new_n840_));
  OR3_X1    g639(.A1(new_n840_), .A2(G113gat), .A3(new_n570_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1340gat));
  OAI21_X1  g641(.A(G120gat), .B1(new_n838_), .B2(new_n280_), .ZN(new_n843_));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n280_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n837_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n844_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(G1341gat));
  OAI21_X1  g646(.A(G127gat), .B1(new_n838_), .B2(new_n622_), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n840_), .A2(G127gat), .A3(new_n622_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1342gat));
  OAI21_X1  g649(.A(G134gat), .B1(new_n838_), .B2(new_n607_), .ZN(new_n851_));
  OR3_X1    g650(.A1(new_n840_), .A2(G134gat), .A3(new_n596_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1343gat));
  NAND4_X1  g652(.A1(new_n507_), .A2(new_n510_), .A3(new_n528_), .A4(new_n505_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n835_), .B2(new_n829_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n717_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n281_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n630_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1346gat));
  AOI21_X1  g661(.A(G162gat), .B1(new_n855_), .B2(new_n603_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n664_), .A2(G162gat), .A3(new_n665_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT122), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n855_), .B2(new_n865_), .ZN(G1347gat));
  NOR3_X1   g665(.A1(new_n440_), .A2(new_n505_), .A3(new_n510_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n717_), .B(new_n867_), .C1(new_n827_), .C2(new_n830_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT62), .B1(new_n868_), .B2(KEYINPUT22), .ZN(new_n869_));
  OAI21_X1  g668(.A(G169gat), .B1(new_n868_), .B2(KEYINPUT62), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT62), .B(G169gat), .C1(new_n868_), .C2(KEYINPUT22), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1348gat));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n874_));
  INV_X1    g673(.A(new_n867_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n835_), .B2(new_n829_), .ZN(new_n876_));
  INV_X1    g675(.A(G176gat), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n280_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n874_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n876_), .A2(new_n874_), .A3(new_n878_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n281_), .B(new_n867_), .C1(new_n827_), .C2(new_n830_), .ZN(new_n881_));
  AOI211_X1 g680(.A(new_n879_), .B(new_n880_), .C1(new_n877_), .C2(new_n881_), .ZN(G1349gat));
  AOI21_X1  g681(.A(G183gat), .B1(new_n876_), .B2(new_n630_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n831_), .A2(new_n875_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n394_), .A2(new_n396_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n630_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n883_), .B1(new_n884_), .B2(new_n887_), .ZN(G1350gat));
  NAND3_X1  g687(.A1(new_n884_), .A2(new_n392_), .A3(new_n603_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n608_), .B(new_n867_), .C1(new_n827_), .C2(new_n830_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n890_), .A2(new_n891_), .A3(G190gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n890_), .B2(G190gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n889_), .B1(new_n892_), .B2(new_n893_), .ZN(G1351gat));
  NAND4_X1  g693(.A1(new_n486_), .A2(new_n511_), .A3(new_n507_), .A4(new_n528_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n835_), .B2(new_n829_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n717_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n281_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT126), .B1(new_n901_), .B2(new_n284_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n630_), .B1(new_n901_), .B2(new_n284_), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT125), .Z(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n896_), .B2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n901_), .A2(new_n284_), .A3(KEYINPUT126), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1354gat));
  NAND2_X1  g706(.A1(new_n896_), .A2(new_n603_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT127), .B(G218gat), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n607_), .A2(new_n909_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n908_), .A2(new_n909_), .B1(new_n896_), .B2(new_n910_), .ZN(G1355gat));
endmodule


