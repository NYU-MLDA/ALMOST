//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT13), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G230gat), .A2(G233gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT64), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT8), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR4_X1   g012(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT66), .A2(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT6), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(KEYINPUT67), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT67), .B1(new_n219_), .B2(new_n221_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n208_), .B(new_n213_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n217_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT7), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n216_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(KEYINPUT68), .A3(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n226_), .A2(new_n232_), .A3(new_n221_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n213_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT8), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n233_), .B2(new_n213_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n224_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G64gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n240_));
  XOR2_X1   g039(.A(G71gat), .B(G78gat), .Z(new_n241_));
  OR2_X1    g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n241_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n212_), .B1(new_n211_), .B2(KEYINPUT9), .ZN(new_n246_));
  INV_X1    g045(.A(new_n211_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT9), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n247_), .A2(KEYINPUT65), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT65), .B1(new_n247_), .B2(new_n248_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n246_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT10), .B(G99gat), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n217_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n221_), .A3(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n238_), .A2(new_n245_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n245_), .B1(new_n238_), .B2(new_n254_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n207_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT70), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n259_), .B(new_n207_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n254_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n233_), .A2(new_n213_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT69), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(KEYINPUT8), .A3(new_n235_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n262_), .B1(new_n265_), .B2(new_n224_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n207_), .B1(new_n266_), .B2(new_n245_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT12), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n238_), .A2(new_n254_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n245_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AOI211_X1 g070(.A(KEYINPUT12), .B(new_n245_), .C1(new_n238_), .C2(new_n254_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n267_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(KEYINPUT71), .B(new_n267_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n261_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G120gat), .B(G148gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G176gat), .B(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n261_), .A2(new_n275_), .A3(new_n276_), .A4(new_n282_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n204_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n277_), .A2(new_n283_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n285_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n291_), .A2(KEYINPUT74), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(KEYINPUT74), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT25), .B(G183gat), .ZN(new_n296_));
  INV_X1    g095(.A(G190gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT26), .B1(new_n297_), .B2(KEYINPUT81), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n297_), .A2(KEYINPUT26), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n296_), .B(new_n298_), .C1(new_n299_), .C2(KEYINPUT81), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(G169gat), .B2(G176gat), .ZN(new_n302_));
  INV_X1    g101(.A(G169gat), .ZN(new_n303_));
  INV_X1    g102(.A(G176gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n307_));
  INV_X1    g106(.A(G183gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT23), .B1(new_n308_), .B2(new_n297_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(G183gat), .A3(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  AND4_X1   g111(.A1(new_n300_), .A2(new_n306_), .A3(new_n307_), .A4(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(KEYINPUT82), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(new_n309_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(G183gat), .B2(G190gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G169gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n313_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT30), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(KEYINPUT84), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT31), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(KEYINPUT84), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G227gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G15gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT83), .B(G43gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G71gat), .B(G99gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT85), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n332_), .B(new_n333_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(KEYINPUT85), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n331_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n331_), .A2(new_n337_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n323_), .A2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n322_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G155gat), .B(G162gat), .Z(new_n344_));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(new_n348_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n346_), .A2(new_n349_), .A3(new_n351_), .A4(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n358_), .B(new_n359_), .C1(new_n350_), .C2(KEYINPUT2), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n344_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n353_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT87), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n337_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n353_), .A2(new_n361_), .A3(new_n336_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT4), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT4), .B1(new_n363_), .B2(new_n337_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G1gat), .B(G29gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n370_), .B1(new_n366_), .B2(KEYINPUT4), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n373_), .B1(new_n383_), .B2(new_n369_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n380_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n343_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n312_), .B1(G183gat), .B2(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n318_), .ZN(new_n390_));
  XOR2_X1   g189(.A(KEYINPUT26), .B(G190gat), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n296_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n315_), .A2(new_n307_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT92), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n305_), .B1(new_n302_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n395_), .B2(new_n302_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n390_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G197gat), .B(G204gat), .Z(new_n399_));
  INV_X1    g198(.A(KEYINPUT90), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT21), .ZN(new_n401_));
  XOR2_X1   g200(.A(G211gat), .B(G218gat), .Z(new_n402_));
  OR2_X1    g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n402_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n399_), .A2(KEYINPUT21), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n388_), .B1(new_n398_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n319_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G226gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT19), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n398_), .A2(new_n406_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n412_), .A2(new_n388_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n414_), .B(new_n415_), .C1(new_n319_), .C2(new_n408_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n413_), .A2(new_n416_), .A3(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n319_), .A2(new_n408_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n398_), .A2(new_n406_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n415_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n412_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n421_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT27), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n398_), .B2(new_n406_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n412_), .B1(new_n435_), .B2(new_n424_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n407_), .A2(new_n409_), .A3(new_n428_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n423_), .B(KEYINPUT27), .C1(new_n438_), .C2(new_n422_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT91), .ZN(new_n441_));
  XOR2_X1   g240(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n442_));
  OR3_X1    g241(.A1(new_n363_), .A2(KEYINPUT29), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n362_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT29), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n442_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G22gat), .B(G50gat), .Z(new_n449_));
  NAND3_X1  g248(.A1(new_n443_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n441_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G228gat), .A2(G233gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n406_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n363_), .A2(KEYINPUT29), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(KEYINPUT89), .ZN(new_n457_));
  OR3_X1    g256(.A1(new_n445_), .A2(KEYINPUT89), .A3(new_n446_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n362_), .A2(KEYINPUT29), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n454_), .B1(new_n406_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G78gat), .B(G106gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n443_), .A2(new_n448_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n449_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT91), .A3(new_n450_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n459_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n453_), .A2(new_n466_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n450_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n464_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n474_));
  AOI211_X1 g273(.A(new_n461_), .B(new_n465_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n473_), .B(new_n441_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n476_));
  AOI211_X1 g275(.A(KEYINPUT98), .B(new_n440_), .C1(new_n472_), .C2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT98), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n476_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n440_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n387_), .B1(new_n477_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT99), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(KEYINPUT99), .B(new_n387_), .C1(new_n477_), .C2(new_n481_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n380_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT33), .B1(new_n384_), .B2(new_n380_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n383_), .A2(new_n369_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n366_), .A2(new_n368_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(new_n381_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n431_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n413_), .A2(new_n416_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT96), .ZN(new_n499_));
  OAI22_X1  g298(.A1(new_n495_), .A2(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n500_), .B1(new_n499_), .B2(new_n498_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n490_), .A2(new_n494_), .B1(new_n386_), .B2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n472_), .A2(new_n476_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT97), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n487_), .B1(new_n375_), .B2(new_n381_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n384_), .A2(KEYINPUT33), .A3(new_n380_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n494_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n498_), .A2(new_n499_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n500_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n375_), .A2(new_n381_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n508_), .B(new_n509_), .C1(new_n510_), .C2(new_n486_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n479_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n386_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n503_), .A2(new_n515_), .A3(new_n480_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n504_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n484_), .A2(new_n485_), .B1(new_n517_), .B2(new_n343_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G29gat), .B(G36gat), .Z(new_n519_));
  XOR2_X1   g318(.A(G43gat), .B(G50gat), .Z(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT15), .Z(new_n522_));
  XOR2_X1   g321(.A(KEYINPUT77), .B(G8gat), .Z(new_n523_));
  INV_X1    g322(.A(G1gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G1gat), .B(G8gat), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n522_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n521_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n532_), .B(new_n535_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G169gat), .B(G197gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n538_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT80), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT80), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n551_), .A3(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n295_), .A2(new_n518_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n269_), .A2(new_n521_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n521_), .B(KEYINPUT15), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n238_), .B2(new_n254_), .ZN(new_n559_));
  OAI211_X1 g358(.A(KEYINPUT35), .B(new_n556_), .C1(new_n557_), .C2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n266_), .A2(new_n535_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .A4(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT76), .Z(new_n571_));
  NAND3_X1  g370(.A1(new_n560_), .A2(new_n565_), .A3(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n560_), .A2(new_n565_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n568_), .B(KEYINPUT36), .Z(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT37), .B(new_n572_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n560_), .A2(new_n565_), .A3(new_n571_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n560_), .B2(new_n565_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n532_), .B(new_n245_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT78), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n581_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585_));
  XOR2_X1   g384(.A(G127gat), .B(G155gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  OR3_X1    g389(.A1(new_n584_), .A2(new_n585_), .A3(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(KEYINPUT17), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n584_), .A2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n580_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n554_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n524_), .A3(new_n386_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n294_), .A2(new_n549_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n577_), .A2(new_n578_), .ZN(new_n603_));
  NOR4_X1   g402(.A1(new_n602_), .A2(new_n518_), .A3(new_n595_), .A4(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n524_), .B1(new_n604_), .B2(new_n386_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n600_), .A2(new_n601_), .A3(new_n605_), .ZN(G1324gat));
  NAND3_X1  g405(.A1(new_n597_), .A2(new_n523_), .A3(new_n440_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n440_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n608_), .A2(new_n609_), .A3(G8gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n608_), .B2(G8gat), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT40), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n607_), .B(KEYINPUT40), .C1(new_n610_), .C2(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1325gat));
  INV_X1    g415(.A(G15gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n343_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n604_), .B2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT41), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n597_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1326gat));
  INV_X1    g421(.A(G22gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n479_), .B(KEYINPUT101), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n597_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n604_), .A2(new_n624_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n627_), .B2(G22gat), .ZN(new_n628_));
  AOI211_X1 g427(.A(KEYINPUT42), .B(new_n623_), .C1(new_n604_), .C2(new_n624_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n625_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(G1327gat));
  INV_X1    g431(.A(new_n603_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n594_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n554_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n386_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n580_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT43), .B1(new_n518_), .B2(new_n638_), .ZN(new_n639_));
  AOI22_X1  g438(.A1(new_n507_), .A2(new_n511_), .B1(new_n476_), .B2(new_n472_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n516_), .B1(new_n640_), .B2(new_n513_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n502_), .A2(KEYINPUT97), .A3(new_n503_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n343_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT98), .B1(new_n503_), .B2(new_n440_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n479_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT99), .B1(new_n646_), .B2(new_n387_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n485_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n643_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n580_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n639_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n294_), .A2(new_n595_), .A3(new_n549_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT44), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  AOI211_X1 g455(.A(new_n656_), .B(new_n653_), .C1(new_n639_), .C2(new_n651_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n386_), .A2(G29gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n637_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  INV_X1    g460(.A(G36gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n658_), .B2(new_n440_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n440_), .A2(KEYINPUT103), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n440_), .A2(KEYINPUT103), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n554_), .A2(new_n662_), .A3(new_n634_), .A4(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n661_), .B1(new_n663_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n668_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n667_), .B(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n655_), .A2(new_n657_), .A3(new_n480_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT46), .B(new_n672_), .C1(new_n673_), .C2(new_n662_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n674_), .ZN(G1329gat));
  INV_X1    g474(.A(G43gat), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n343_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n658_), .A2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n635_), .B2(new_n343_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n678_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1330gat));
  AOI21_X1  g484(.A(G50gat), .B1(new_n636_), .B2(new_n624_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n503_), .A2(G50gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n658_), .B2(new_n687_), .ZN(G1331gat));
  INV_X1    g487(.A(new_n553_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n294_), .A2(new_n595_), .A3(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(new_n633_), .A3(new_n649_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT109), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(KEYINPUT109), .ZN(new_n693_));
  INV_X1    g492(.A(G57gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n515_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n692_), .A2(new_n693_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n691_), .B(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(KEYINPUT110), .A3(new_n695_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n518_), .B2(new_n549_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n549_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n649_), .A2(KEYINPUT106), .A3(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n704_), .A2(new_n706_), .A3(new_n596_), .A4(new_n295_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n515_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n649_), .A2(new_n705_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n294_), .B1(new_n710_), .B2(new_n703_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n711_), .A2(KEYINPUT107), .A3(new_n596_), .A4(new_n706_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT108), .B1(new_n713_), .B2(new_n694_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n715_), .B(G57gat), .C1(new_n709_), .C2(new_n712_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n702_), .A2(new_n714_), .A3(new_n716_), .ZN(G1332gat));
  INV_X1    g516(.A(new_n707_), .ZN(new_n718_));
  INV_X1    g517(.A(G64gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n666_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n700_), .A2(new_n666_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(G64gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT48), .B(new_n719_), .C1(new_n700_), .C2(new_n666_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(G1333gat));
  INV_X1    g524(.A(G71gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n718_), .A2(new_n726_), .A3(new_n618_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT49), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n700_), .A2(new_n618_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G71gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT49), .B(new_n726_), .C1(new_n700_), .C2(new_n618_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n700_), .A2(new_n624_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n733_), .A2(G78gat), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n733_), .B2(G78gat), .ZN(new_n736_));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n624_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT112), .ZN(new_n739_));
  OAI22_X1  g538(.A1(new_n735_), .A2(new_n736_), .B1(new_n707_), .B2(new_n739_), .ZN(G1335gat));
  AND2_X1   g539(.A1(new_n711_), .A2(new_n706_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n634_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n386_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n294_), .A2(new_n594_), .A3(new_n549_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n652_), .A2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT113), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n515_), .A2(new_n209_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1336gat));
  AOI21_X1  g548(.A(G92gat), .B1(new_n743_), .B2(new_n440_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n666_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(new_n210_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n747_), .B2(new_n752_), .ZN(G1337gat));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n755_));
  OAI21_X1  g554(.A(G99gat), .B1(new_n746_), .B2(new_n343_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n618_), .A2(new_n252_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n711_), .A2(new_n634_), .A3(new_n706_), .A4(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n755_), .B1(new_n756_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT115), .Z(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n760_), .B(new_n763_), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n652_), .A2(new_n503_), .A3(new_n745_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(G106gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G106gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n503_), .A2(new_n217_), .ZN(new_n769_));
  OAI22_X1  g568(.A1(new_n767_), .A2(new_n768_), .B1(new_n742_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  OAI221_X1 g571(.A(new_n772_), .B1(new_n742_), .B2(new_n769_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT119), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n689_), .A2(G113gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n646_), .A2(new_n618_), .A3(new_n386_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n275_), .A2(new_n778_), .A3(new_n276_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n238_), .A2(new_n245_), .A3(new_n254_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n206_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT12), .B1(new_n266_), .B2(new_n245_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n269_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n207_), .A2(new_n781_), .B1(new_n785_), .B2(KEYINPUT55), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n779_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n283_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  AOI211_X1 g588(.A(new_n789_), .B(new_n282_), .C1(new_n779_), .C2(new_n786_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n534_), .A2(new_n536_), .A3(new_n540_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n545_), .B1(new_n539_), .B2(new_n537_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n548_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n285_), .A2(new_n791_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n791_), .B1(new_n285_), .B2(new_n795_), .ZN(new_n798_));
  OAI22_X1  g597(.A1(new_n788_), .A2(new_n790_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n580_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n787_), .A2(new_n283_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n789_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n283_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n798_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n796_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT58), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n285_), .A2(new_n549_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n795_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n288_), .B2(new_n285_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n603_), .B1(new_n811_), .B2(new_n814_), .ZN(new_n815_));
  OAI22_X1  g614(.A1(new_n801_), .A2(new_n808_), .B1(new_n815_), .B2(KEYINPUT57), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n809_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n633_), .B1(new_n817_), .B2(new_n813_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n595_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n575_), .A2(new_n553_), .A3(new_n579_), .A4(new_n594_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n290_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n288_), .A2(new_n285_), .B1(new_n202_), .B2(new_n203_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT116), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n291_), .A2(new_n828_), .A3(new_n823_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n827_), .A2(new_n829_), .A3(KEYINPUT54), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT54), .B1(new_n827_), .B2(new_n829_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI211_X1 g631(.A(KEYINPUT59), .B(new_n777_), .C1(new_n821_), .C2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n777_), .B1(new_n821_), .B2(new_n832_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n828_), .B1(new_n291_), .B2(new_n823_), .ZN(new_n839_));
  AOI211_X1 g638(.A(KEYINPUT116), .B(new_n822_), .C1(new_n287_), .C2(new_n290_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n827_), .A2(new_n829_), .A3(KEYINPUT54), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n818_), .A2(new_n819_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n815_), .A2(KEYINPUT57), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n799_), .A2(new_n800_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n805_), .A2(new_n807_), .A3(KEYINPUT58), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n580_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n844_), .A2(new_n845_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n843_), .B1(new_n595_), .B2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n850_), .C2(new_n777_), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n776_), .B(new_n833_), .C1(new_n837_), .C2(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n850_), .A2(new_n705_), .A3(new_n777_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(G113gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n775_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n854_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n837_), .A2(new_n851_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n821_), .A2(new_n832_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n777_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n836_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT119), .B(new_n856_), .C1(new_n861_), .C2(new_n776_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n855_), .A2(new_n862_), .ZN(G1340gat));
  INV_X1    g662(.A(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n294_), .B2(KEYINPUT60), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n835_), .B(new_n865_), .C1(KEYINPUT60), .C2(new_n864_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n860_), .A2(new_n295_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n837_), .B2(new_n851_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869_));
  OAI21_X1  g668(.A(G120gat), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  AOI211_X1 g669(.A(KEYINPUT120), .B(new_n867_), .C1(new_n837_), .C2(new_n851_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n866_), .B1(new_n870_), .B2(new_n871_), .ZN(G1341gat));
  OAI21_X1  g671(.A(G127gat), .B1(new_n861_), .B2(new_n595_), .ZN(new_n873_));
  INV_X1    g672(.A(G127gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n835_), .A2(new_n874_), .A3(new_n594_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1342gat));
  XOR2_X1   g675(.A(KEYINPUT121), .B(G134gat), .Z(new_n877_));
  NOR3_X1   g676(.A1(new_n861_), .A2(new_n638_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G134gat), .B1(new_n835_), .B2(new_n603_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n618_), .A2(new_n479_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n858_), .A2(new_n386_), .A3(new_n751_), .A4(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n705_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT122), .B(G141gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1344gat));
  NOR2_X1   g684(.A1(new_n882_), .A2(new_n294_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n348_), .ZN(G1345gat));
  OR3_X1    g686(.A1(new_n882_), .A2(KEYINPUT123), .A3(new_n595_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT123), .B1(new_n882_), .B2(new_n595_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT124), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n890_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n888_), .A2(new_n889_), .A3(new_n892_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1346gat));
  OAI21_X1  g695(.A(G162gat), .B1(new_n882_), .B2(new_n638_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n633_), .A2(G162gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n882_), .B2(new_n898_), .ZN(G1347gat));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n387_), .A2(new_n666_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT125), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n624_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n858_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n705_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT22), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n900_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G169gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n303_), .B1(new_n905_), .B2(new_n900_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n907_), .B2(new_n909_), .ZN(G1348gat));
  INV_X1    g709(.A(new_n904_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n304_), .A3(new_n295_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n858_), .A2(new_n479_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n913_), .A2(new_n294_), .A3(new_n902_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n914_), .B2(new_n304_), .ZN(G1349gat));
  NOR3_X1   g714(.A1(new_n904_), .A2(new_n595_), .A3(new_n296_), .ZN(new_n916_));
  OR3_X1    g715(.A1(new_n913_), .A2(new_n595_), .A3(new_n902_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n308_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n904_), .B2(new_n638_), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT126), .Z(new_n920_));
  NAND3_X1  g719(.A1(new_n911_), .A2(new_n603_), .A3(new_n392_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1351gat));
  AND2_X1   g721(.A1(new_n858_), .A2(new_n881_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n751_), .A2(new_n386_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n549_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n295_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g729(.A(KEYINPUT63), .B(G211gat), .C1(new_n926_), .C2(new_n594_), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT63), .B(G211gat), .Z(new_n932_));
  AND3_X1   g731(.A1(new_n926_), .A2(new_n594_), .A3(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1354gat));
  AND3_X1   g733(.A1(new_n926_), .A2(G218gat), .A3(new_n580_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n925_), .A2(KEYINPUT127), .A3(new_n633_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(G218gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT127), .B1(new_n925_), .B2(new_n633_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n935_), .B1(new_n937_), .B2(new_n938_), .ZN(G1355gat));
endmodule


