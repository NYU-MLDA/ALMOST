//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(KEYINPUT77), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  INV_X1    g012(.A(G1gat), .ZN(new_n214_));
  INV_X1    g013(.A(G8gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(KEYINPUT77), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n218_), .B1(new_n212_), .B2(new_n219_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n210_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT15), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n210_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(new_n219_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n217_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n208_), .A2(KEYINPUT15), .A3(new_n209_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n220_), .A4(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n223_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n210_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n227_), .A2(new_n232_), .A3(new_n220_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n230_), .B1(new_n223_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n205_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n223_), .A2(new_n233_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n230_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n223_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n204_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n235_), .A2(KEYINPUT80), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT80), .B1(new_n235_), .B2(new_n240_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G230gat), .A2(G233gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT6), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT6), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(G99gat), .A3(G106gat), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT65), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT65), .B1(new_n246_), .B2(new_n248_), .ZN(new_n250_));
  AND2_X1   g049(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n251_), .A2(new_n252_), .A3(G106gat), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n249_), .A2(new_n250_), .A3(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G85gat), .A2(G92gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G85gat), .A2(G92gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n257_), .B2(KEYINPUT9), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT9), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n259_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n256_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n258_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n254_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n257_), .A2(new_n255_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT8), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n249_), .A2(new_n250_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT7), .ZN(new_n269_));
  INV_X1    g068(.A(G99gat), .ZN(new_n270_));
  INV_X1    g069(.A(G106gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n267_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n247_), .B1(G99gat), .B2(G106gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n245_), .A2(KEYINPUT6), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n272_), .B(new_n273_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n266_), .B1(new_n278_), .B2(new_n265_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n264_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G57gat), .B(G64gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G71gat), .B(G78gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT11), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(KEYINPUT11), .B2(new_n281_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n281_), .A2(KEYINPUT11), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n284_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT66), .B1(new_n280_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n285_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n283_), .B1(new_n290_), .B2(new_n286_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n291_), .B(new_n264_), .C1(new_n275_), .C2(new_n279_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n244_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n292_), .B2(new_n289_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n292_), .A2(new_n244_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT12), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n280_), .B2(new_n288_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT65), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT65), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n274_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n267_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n246_), .A2(new_n248_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n272_), .A2(new_n273_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n265_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT8), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n303_), .A2(new_n307_), .B1(new_n263_), .B2(new_n254_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n308_), .A2(KEYINPUT12), .A3(new_n291_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n295_), .B1(new_n297_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n294_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G120gat), .B(G148gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G176gat), .B(G204gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT68), .Z(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n294_), .A2(new_n316_), .A3(new_n310_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n323_));
  OAI22_X1  g122(.A1(new_n322_), .A2(new_n323_), .B1(KEYINPUT70), .B2(KEYINPUT13), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n321_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G15gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G71gat), .B(G99gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT84), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT22), .B(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT83), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n338_), .A2(KEYINPUT83), .A3(new_n339_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT23), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(G183gat), .B2(G190gat), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n342_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT25), .B(G183gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G190gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n351_));
  INV_X1    g150(.A(G169gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n337_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n339_), .A2(KEYINPUT24), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n350_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n345_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT24), .B1(new_n353_), .B2(new_n354_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n344_), .B(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT82), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n357_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n335_), .B1(new_n347_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n365_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n357_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n342_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(KEYINPUT84), .A3(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n367_), .A2(new_n372_), .A3(KEYINPUT30), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT30), .B1(new_n367_), .B2(new_n372_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT85), .B(G43gat), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n347_), .A2(new_n335_), .A3(new_n366_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT84), .B1(new_n370_), .B2(new_n371_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n367_), .A2(new_n372_), .A3(KEYINPUT30), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n377_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n334_), .B1(new_n376_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n375_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n382_), .A3(new_n377_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n333_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT86), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G127gat), .B(G134gat), .Z(new_n389_));
  XOR2_X1   g188(.A(G113gat), .B(G120gat), .Z(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT31), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n384_), .A2(KEYINPUT86), .A3(new_n387_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n392_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n396_), .B2(new_n388_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT87), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G57gat), .B(G85gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(G141gat), .ZN(new_n406_));
  INV_X1    g205(.A(G148gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT3), .ZN(new_n409_));
  OR3_X1    g208(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT2), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n409_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(KEYINPUT88), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G155gat), .B(G162gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n389_), .B(new_n390_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n418_), .A2(KEYINPUT1), .ZN(new_n422_));
  NAND3_X1  g221(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n408_), .A2(new_n423_), .A3(new_n411_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n420_), .A2(new_n421_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n418_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n391_), .B1(new_n428_), .B2(new_n425_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n429_), .A3(KEYINPUT4), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n420_), .A2(new_n426_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n391_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n405_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n427_), .A2(new_n429_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n405_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n404_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT96), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT33), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n404_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n430_), .A2(new_n433_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n436_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G226gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT19), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n349_), .B(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n348_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT93), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n355_), .B1(new_n453_), .B2(new_n356_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n453_), .B2(new_n356_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n359_), .A2(new_n345_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT94), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT94), .B1(new_n359_), .B2(new_n345_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n452_), .B(new_n455_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n340_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n346_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G211gat), .B(G218gat), .Z(new_n464_));
  INV_X1    g263(.A(KEYINPUT21), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G197gat), .B(G204gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G204gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(G197gat), .B(G204gat), .Z(new_n470_));
  OAI211_X1 g269(.A(KEYINPUT21), .B(new_n469_), .C1(new_n470_), .C2(KEYINPUT89), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n464_), .A3(KEYINPUT21), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT20), .B1(new_n463_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n474_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n449_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT18), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G64gat), .B(G92gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n463_), .B2(new_n474_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n367_), .A2(new_n372_), .A3(new_n476_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n448_), .A3(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n478_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n483_), .B1(new_n478_), .B2(new_n487_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n474_), .A2(KEYINPUT90), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n472_), .A2(new_n492_), .A3(new_n473_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT20), .B1(new_n463_), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n448_), .B1(new_n495_), .B2(new_n477_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n485_), .A2(new_n449_), .A3(new_n486_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n482_), .A2(KEYINPUT32), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n443_), .A2(new_n436_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n501_), .B(new_n403_), .C1(new_n436_), .C2(new_n435_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n498_), .A2(new_n500_), .B1(new_n502_), .B2(new_n438_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n460_), .A2(new_n462_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n484_), .B1(new_n504_), .B2(new_n476_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n474_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n448_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n485_), .A2(new_n448_), .A3(new_n486_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n499_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n446_), .A2(new_n490_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(G228gat), .ZN(new_n511_));
  INV_X1    g310(.A(G233gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n476_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n431_), .A2(KEYINPUT29), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n491_), .A2(new_n493_), .B1(new_n431_), .B2(KEYINPUT29), .ZN(new_n517_));
  INV_X1    g316(.A(new_n513_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G22gat), .B(G50gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n516_), .B(new_n522_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  OR4_X1    g323(.A1(KEYINPUT28), .A2(new_n428_), .A3(KEYINPUT29), .A4(new_n425_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT28), .B1(new_n431_), .B2(KEYINPUT29), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G78gat), .B(G106gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT91), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n524_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n521_), .A2(new_n531_), .A3(new_n523_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n498_), .A2(new_n483_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n482_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT27), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT27), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n502_), .A2(new_n438_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n535_), .A2(new_n543_), .ZN(new_n544_));
  OAI22_X1  g343(.A1(new_n510_), .A2(new_n535_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT87), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n394_), .B(new_n546_), .C1(new_n396_), .C2(new_n388_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n398_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT97), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n541_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n538_), .A2(new_n540_), .A3(KEYINPUT97), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n397_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n535_), .A2(new_n542_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI211_X1 g354(.A(new_n243_), .B(new_n329_), .C1(new_n548_), .C2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  OAI22_X1  g358(.A1(new_n280_), .A2(new_n232_), .B1(KEYINPUT35), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT72), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT72), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n280_), .A2(new_n228_), .A3(new_n225_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT74), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n567_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n570_), .B2(new_n560_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n561_), .A2(KEYINPUT74), .A3(new_n567_), .A4(new_n565_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n566_), .A2(new_n568_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT73), .ZN(new_n575_));
  XOR2_X1   g374(.A(G134gat), .B(G162gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(KEYINPUT36), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n577_), .B(KEYINPUT36), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n573_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT37), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  INV_X1    g383(.A(new_n581_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT75), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n585_), .B1(new_n573_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n566_), .A2(new_n568_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n572_), .A2(new_n571_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n588_), .A2(new_n586_), .A3(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n584_), .B(new_n579_), .C1(new_n587_), .C2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT76), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n583_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n583_), .B2(new_n591_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n227_), .A2(new_n220_), .ZN(new_n596_));
  INV_X1    g395(.A(G231gat), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(new_n512_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n288_), .A2(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n599_), .B(new_n283_), .C1(new_n290_), .C2(new_n286_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n596_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT78), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n291_), .A2(new_n598_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(new_n220_), .A3(new_n227_), .A4(new_n601_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n608_));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT16), .ZN(new_n610_));
  XOR2_X1   g409(.A(G183gat), .B(G211gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n607_), .A2(new_n608_), .A3(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n607_), .A2(new_n612_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n603_), .A2(new_n606_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT17), .B1(new_n615_), .B2(new_n612_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n613_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT79), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT79), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n619_), .B(new_n613_), .C1(new_n614_), .C2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n595_), .A2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n556_), .A2(new_n622_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n623_), .A2(KEYINPUT98), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(KEYINPUT98), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n624_), .A2(new_n214_), .A3(new_n542_), .A4(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n548_), .A2(new_n555_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n587_), .A2(new_n590_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(new_n579_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n629_), .A2(KEYINPUT99), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT99), .B1(new_n629_), .B2(new_n632_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n235_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n240_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n329_), .A2(new_n621_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n543_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n626_), .A2(new_n627_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n628_), .A2(new_n641_), .A3(new_n642_), .ZN(G1324gat));
  INV_X1    g442(.A(new_n552_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n644_), .B(new_n639_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT100), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(G8gat), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT39), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n647_), .A2(new_n651_), .A3(G8gat), .A4(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n624_), .A2(new_n215_), .A3(new_n644_), .A4(new_n625_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(KEYINPUT40), .A3(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1325gat));
  NAND2_X1  g458(.A1(new_n398_), .A2(new_n547_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G15gat), .B1(new_n640_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT41), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n624_), .A2(new_n625_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n664_), .A2(G15gat), .A3(new_n661_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n663_), .A2(new_n665_), .ZN(G1326gat));
  INV_X1    g465(.A(new_n535_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G22gat), .B1(new_n640_), .B2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(KEYINPUT42), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(KEYINPUT42), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n667_), .A2(G22gat), .ZN(new_n671_));
  OAI22_X1  g470(.A1(new_n669_), .A2(new_n670_), .B1(new_n664_), .B2(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(new_n621_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n632_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n556_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n542_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n329_), .A2(new_n673_), .A3(new_n638_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n629_), .A2(new_n679_), .A3(new_n595_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n629_), .B2(new_n595_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT44), .B(new_n678_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n542_), .A2(G29gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n677_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  NOR3_X1   g487(.A1(new_n675_), .A2(G36gat), .A3(new_n552_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n684_), .A2(new_n644_), .A3(new_n685_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n692_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT101), .B1(new_n692_), .B2(G36gat), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT103), .B(new_n691_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT103), .B1(new_n698_), .B2(KEYINPUT104), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n697_), .A2(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(G1329gat));
  NAND3_X1  g500(.A1(new_n686_), .A2(G43gat), .A3(new_n553_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT105), .B(G43gat), .Z(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n675_), .B2(new_n661_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g505(.A1(new_n675_), .A2(G50gat), .A3(new_n667_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n686_), .A2(new_n535_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G50gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G50gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1331gat));
  NAND4_X1  g511(.A1(new_n635_), .A2(new_n673_), .A3(new_n329_), .A4(new_n243_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n543_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n629_), .A2(new_n638_), .ZN(new_n715_));
  NOR4_X1   g514(.A1(new_n715_), .A2(new_n621_), .A3(new_n595_), .A4(new_n328_), .ZN(new_n716_));
  INV_X1    g515(.A(G57gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n542_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n718_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n713_), .B2(new_n552_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT48), .ZN(new_n721_));
  INV_X1    g520(.A(G64gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n716_), .A2(new_n722_), .A3(new_n644_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n713_), .B2(new_n661_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT49), .ZN(new_n726_));
  INV_X1    g525(.A(G71gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n716_), .A2(new_n727_), .A3(new_n660_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1334gat));
  OAI21_X1  g528(.A(G78gat), .B1(new_n713_), .B2(new_n667_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT50), .ZN(new_n731_));
  INV_X1    g530(.A(G78gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n716_), .A2(new_n732_), .A3(new_n535_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1335gat));
  OR2_X1    g533(.A1(new_n680_), .A2(new_n681_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n638_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n328_), .A2(new_n673_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n543_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n629_), .A2(new_n329_), .A3(new_n638_), .A4(new_n674_), .ZN(new_n740_));
  OR3_X1    g539(.A1(new_n740_), .A2(G85gat), .A3(new_n543_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1336gat));
  OAI21_X1  g541(.A(G92gat), .B1(new_n738_), .B2(new_n552_), .ZN(new_n743_));
  OR3_X1    g542(.A1(new_n740_), .A2(G92gat), .A3(new_n552_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n738_), .B2(new_n661_), .ZN(new_n746_));
  OR3_X1    g545(.A1(new_n397_), .A2(new_n252_), .A3(new_n251_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n740_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(KEYINPUT107), .A2(KEYINPUT51), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n748_), .B(new_n749_), .Z(G1338gat));
  OAI21_X1  g549(.A(G106gat), .B1(new_n738_), .B2(new_n667_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT52), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(KEYINPUT52), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n535_), .A2(new_n271_), .ZN(new_n754_));
  OAI22_X1  g553(.A1(new_n752_), .A2(new_n753_), .B1(new_n740_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g555(.A(KEYINPUT59), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n618_), .A2(new_n243_), .A3(new_n620_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n618_), .A2(new_n243_), .A3(KEYINPUT108), .A4(new_n620_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n764_));
  XOR2_X1   g563(.A(KEYINPUT109), .B(KEYINPUT54), .Z(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n763_), .B(new_n765_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n631_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n223_), .A2(new_n229_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n230_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n773_), .B2(new_n772_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n204_), .B1(new_n236_), .B2(new_n230_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n637_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n325_), .B2(new_n321_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n736_), .A2(new_n320_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n292_), .A2(new_n244_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT12), .B1(new_n308_), .B2(new_n291_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n301_), .A2(new_n302_), .B1(new_n306_), .B2(KEYINPUT8), .ZN(new_n784_));
  INV_X1    g583(.A(new_n253_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n268_), .A2(new_n263_), .A3(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n296_), .B(new_n288_), .C1(new_n784_), .C2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n782_), .B1(new_n783_), .B2(new_n787_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n784_), .A2(new_n786_), .A3(new_n288_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n783_), .B2(new_n787_), .ZN(new_n790_));
  OAI22_X1  g589(.A1(new_n788_), .A2(KEYINPUT55), .B1(new_n790_), .B2(new_n244_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n310_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n317_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(KEYINPUT110), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT110), .B1(new_n794_), .B2(new_n795_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT56), .B(new_n317_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n310_), .A2(new_n792_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n788_), .A2(KEYINPUT55), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n802_), .B(new_n803_), .C1(new_n244_), .C2(new_n790_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n804_), .A2(KEYINPUT111), .A3(KEYINPUT56), .A4(new_n317_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n801_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n781_), .B1(new_n798_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n780_), .B1(new_n807_), .B2(KEYINPUT112), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n794_), .A2(new_n795_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n794_), .A2(KEYINPUT110), .A3(new_n795_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n801_), .A4(new_n805_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n781_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n771_), .B1(new_n808_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n809_), .A2(new_n819_), .A3(new_n799_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n804_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n317_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n320_), .A3(new_n777_), .A4(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n595_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n779_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n807_), .A2(KEYINPUT112), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n631_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n818_), .B(new_n824_), .C1(new_n827_), .C2(KEYINPUT57), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n769_), .B1(new_n828_), .B2(new_n621_), .ZN(new_n829_));
  NOR4_X1   g628(.A1(new_n644_), .A2(new_n397_), .A3(new_n535_), .A4(new_n543_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n757_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n825_), .A2(new_n826_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n834_), .A2(new_n771_), .B1(new_n595_), .B2(new_n823_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n632_), .B1(new_n808_), .B2(new_n817_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n770_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n673_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT59), .B(new_n830_), .C1(new_n838_), .C2(new_n769_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n833_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(G113gat), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n243_), .ZN(new_n843_));
  OR3_X1    g642(.A1(new_n829_), .A2(KEYINPUT115), .A3(new_n831_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT115), .B1(new_n829_), .B2(new_n831_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n736_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n842_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(KEYINPUT116), .A3(new_n842_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n843_), .B1(new_n849_), .B2(new_n850_), .ZN(G1340gat));
  NOR2_X1   g650(.A1(new_n328_), .A2(KEYINPUT60), .ZN(new_n852_));
  MUX2_X1   g651(.A(new_n852_), .B(KEYINPUT60), .S(G120gat), .Z(new_n853_));
  NAND3_X1  g652(.A1(new_n844_), .A2(new_n845_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n328_), .B1(new_n832_), .B2(new_n839_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G120gat), .B1(new_n855_), .B2(KEYINPUT117), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n857_), .B(new_n328_), .C1(new_n832_), .C2(new_n839_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT118), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n861_), .B(new_n854_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1341gat));
  OAI21_X1  g662(.A(G127gat), .B1(new_n841_), .B2(new_n621_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n621_), .A2(G127gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n844_), .A2(new_n845_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1342gat));
  NAND3_X1  g666(.A1(new_n844_), .A2(new_n631_), .A3(new_n845_), .ZN(new_n868_));
  INV_X1    g667(.A(G134gat), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT119), .B(G134gat), .Z(new_n871_));
  OAI211_X1 g670(.A(new_n595_), .B(new_n871_), .C1(new_n833_), .C2(new_n840_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT120), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n870_), .A2(new_n875_), .A3(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1343gat));
  INV_X1    g676(.A(new_n829_), .ZN(new_n878_));
  NOR4_X1   g677(.A1(new_n660_), .A2(new_n644_), .A3(new_n667_), .A4(new_n543_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n638_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n406_), .ZN(G1344gat));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n328_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n407_), .ZN(G1345gat));
  NOR2_X1   g683(.A1(new_n880_), .A2(new_n621_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT61), .B(G155gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  INV_X1    g686(.A(new_n595_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G162gat), .B1(new_n880_), .B2(new_n888_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n632_), .A2(G162gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n880_), .B2(new_n890_), .ZN(G1347gat));
  AND4_X1   g690(.A1(new_n660_), .A2(new_n878_), .A3(new_n554_), .A4(new_n644_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n352_), .B1(new_n892_), .B2(new_n736_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n893_), .A2(KEYINPUT62), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n336_), .A3(new_n736_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(KEYINPUT62), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(G1348gat));
  AOI22_X1  g696(.A1(new_n892_), .A2(new_n329_), .B1(KEYINPUT121), .B2(G176gat), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT121), .A2(G176gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT122), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n898_), .B(new_n900_), .ZN(G1349gat));
  NAND2_X1  g700(.A1(new_n892_), .A2(new_n673_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(KEYINPUT123), .B2(G183gat), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n348_), .B1(new_n904_), .B2(G183gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n902_), .B2(new_n905_), .ZN(G1350gat));
  NAND2_X1  g705(.A1(new_n892_), .A2(new_n595_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G190gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n892_), .A2(new_n631_), .A3(new_n451_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1351gat));
  XNOR2_X1  g709(.A(KEYINPUT125), .B(G197gat), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n660_), .A2(new_n667_), .A3(new_n542_), .A4(new_n552_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n878_), .A2(new_n912_), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT124), .Z(new_n914_));
  AOI21_X1  g713(.A(new_n911_), .B1(new_n914_), .B2(new_n736_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n913_), .B(KEYINPUT124), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(G197gat), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n916_), .A2(new_n638_), .A3(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n915_), .A2(new_n919_), .ZN(G1352gat));
  NOR2_X1   g719(.A1(new_n916_), .A2(new_n328_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT126), .B(G204gat), .Z(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n921_), .B2(new_n924_), .ZN(G1353gat));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT127), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n621_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n914_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n914_), .B2(new_n928_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1354gat));
  OR3_X1    g730(.A1(new_n916_), .A2(G218gat), .A3(new_n632_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G218gat), .B1(new_n916_), .B2(new_n888_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1355gat));
endmodule


