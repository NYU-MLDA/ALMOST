//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT34), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT35), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT71), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G29gat), .B(G36gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT15), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n216_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n217_), .B(new_n218_), .C1(new_n216_), .C2(KEYINPUT9), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n218_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n224_), .A2(new_n226_), .A3(new_n216_), .A4(KEYINPUT9), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n215_), .A2(new_n219_), .A3(new_n223_), .A4(new_n227_), .ZN(new_n228_));
  OR3_X1    g027(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n229_), .B(new_n230_), .C1(new_n212_), .C2(new_n214_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n218_), .A2(new_n225_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT8), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n231_), .A2(new_n234_), .A3(new_n232_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n233_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n231_), .A2(new_n232_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n228_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n206_), .B1(new_n210_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n209_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(new_n239_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT72), .B1(new_n210_), .B2(new_n239_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n203_), .A2(new_n204_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  OAI221_X1 g046(.A(new_n240_), .B1(new_n241_), .B2(new_n239_), .C1(new_n243_), .C2(new_n245_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G190gat), .B(G218gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT73), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G134gat), .B(G162gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT36), .Z(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n253_), .A2(KEYINPUT36), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n247_), .A2(new_n248_), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(KEYINPUT37), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT74), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n249_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT74), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n254_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n257_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT37), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n259_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G15gat), .B(G22gat), .ZN(new_n268_));
  INV_X1    g067(.A(G1gat), .ZN(new_n269_));
  INV_X1    g068(.A(G8gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT14), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n268_), .B1(new_n271_), .B2(KEYINPUT75), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(KEYINPUT75), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G1gat), .B(G8gat), .ZN(new_n274_));
  OR3_X1    g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n274_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(G231gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT76), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT76), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G71gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G78gat), .ZN(new_n284_));
  INV_X1    g083(.A(G78gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G71gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G57gat), .B(G64gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(KEYINPUT11), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(new_n288_), .B2(KEYINPUT11), .ZN(new_n291_));
  INV_X1    g090(.A(G64gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G57gat), .ZN(new_n293_));
  INV_X1    g092(.A(G57gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G64gat), .ZN(new_n295_));
  AND4_X1   g094(.A1(new_n290_), .A2(new_n293_), .A3(new_n295_), .A4(KEYINPUT11), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n289_), .B1(new_n291_), .B2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n295_), .A3(KEYINPUT11), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT67), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n293_), .A2(new_n295_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT11), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n293_), .A2(new_n295_), .A3(new_n290_), .A4(KEYINPUT11), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n299_), .A2(new_n302_), .A3(new_n287_), .A4(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n297_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n282_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n280_), .A2(new_n281_), .A3(new_n305_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G127gat), .B(G155gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G183gat), .B(G211gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .A4(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n279_), .A2(KEYINPUT79), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n279_), .A2(KEYINPUT79), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n297_), .A2(new_n304_), .A3(KEYINPUT68), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT68), .B1(new_n297_), .B2(new_n304_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n316_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n314_), .B(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n323_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n315_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n267_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n239_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT12), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n320_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n231_), .A2(new_n232_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n234_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n231_), .A2(new_n234_), .A3(new_n232_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n297_), .A2(new_n304_), .A3(KEYINPUT68), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n334_), .A2(new_n339_), .A3(new_n228_), .A4(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G230gat), .A2(G233gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT64), .Z(new_n343_));
  NAND3_X1  g142(.A1(new_n239_), .A2(KEYINPUT12), .A3(new_n306_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n333_), .A2(new_n341_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n343_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n334_), .A2(new_n340_), .B1(new_n339_), .B2(new_n228_), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n239_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G120gat), .B(G148gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT5), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G176gat), .B(G204gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n345_), .A2(new_n349_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT69), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n345_), .A2(new_n349_), .A3(new_n356_), .A4(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n353_), .B1(new_n345_), .B2(new_n349_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT70), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n363_), .A3(new_n360_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(KEYINPUT13), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT13), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n363_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n367_));
  AOI211_X1 g166(.A(KEYINPUT70), .B(new_n359_), .C1(new_n355_), .C2(new_n357_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n330_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G204gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G197gat), .ZN(new_n373_));
  INV_X1    g172(.A(G197gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G204gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G218gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G211gat), .ZN(new_n378_));
  INV_X1    g177(.A(G211gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G218gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n381_), .A3(KEYINPUT21), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n372_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT21), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G197gat), .B(G204gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G211gat), .B(G218gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n376_), .B2(KEYINPUT21), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n382_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT87), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n397_), .A2(KEYINPUT87), .A3(new_n398_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n393_), .B(new_n396_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n402_), .A2(G155gat), .A3(G162gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(G155gat), .B2(G162gat), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n404_), .A2(new_n405_), .B1(G155gat), .B2(G162gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n407_), .A2(KEYINPUT1), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(KEYINPUT1), .ZN(new_n409_));
  INV_X1    g208(.A(new_n405_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n408_), .B(new_n409_), .C1(new_n410_), .C2(new_n403_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n394_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n412_), .A2(new_n397_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n401_), .A2(new_n406_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n390_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n390_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  OAI221_X1 g220(.A(new_n390_), .B1(new_n419_), .B2(new_n418_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n421_), .A2(new_n422_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n414_), .A2(new_n415_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G22gat), .B(G50gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT28), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n429_), .B(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n426_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n432_), .B1(new_n433_), .B2(KEYINPUT90), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n428_), .A2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n425_), .A2(KEYINPUT90), .A3(new_n427_), .A4(new_n432_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n438_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT92), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT21), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n381_), .B1(new_n443_), .B2(new_n386_), .ZN(new_n444_));
  OAI211_X1 g243(.A(KEYINPUT21), .B(new_n383_), .C1(new_n376_), .C2(KEYINPUT88), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n386_), .A2(new_n443_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n444_), .A2(new_n445_), .B1(new_n381_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT25), .B(G183gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT26), .B(G190gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G169gat), .A2(G176gat), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n448_), .A2(new_n449_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n454_));
  AND3_X1   g253(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n456_), .ZN(new_n458_));
  INV_X1    g257(.A(G183gat), .ZN(new_n459_));
  INV_X1    g258(.A(G190gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT22), .ZN(new_n464_));
  INV_X1    g263(.A(G176gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(G169gat), .ZN(new_n466_));
  INV_X1    g265(.A(G169gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n453_), .A2(new_n457_), .B1(new_n463_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT20), .B1(new_n447_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n463_), .A2(new_n469_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT26), .ZN(new_n474_));
  NAND2_X1  g273(.A1(KEYINPUT83), .A2(G183gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT25), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT26), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT25), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(KEYINPUT83), .A3(G183gat), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n474_), .A2(new_n476_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n457_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n452_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT85), .B1(new_n483_), .B2(new_n450_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n467_), .A2(new_n465_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT24), .A4(new_n452_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n472_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(new_n390_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n442_), .B1(new_n471_), .B2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G8gat), .B(G36gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT18), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G64gat), .B(G92gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n438_), .B(new_n439_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT20), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n497_), .B1(new_n447_), .B2(new_n470_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n489_), .A2(new_n390_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n491_), .A2(new_n495_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT93), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n459_), .A2(KEYINPUT25), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n479_), .A2(G183gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n460_), .A2(KEYINPUT26), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n477_), .A2(G190gat), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n455_), .A2(new_n456_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n454_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n485_), .A2(KEYINPUT24), .A3(new_n452_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .A4(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n472_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n390_), .A2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n457_), .A2(new_n481_), .A3(new_n484_), .A4(new_n487_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n386_), .A2(new_n443_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n373_), .A2(new_n375_), .A3(new_n385_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n515_), .B(new_n388_), .C1(new_n516_), .C2(new_n384_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n514_), .A2(new_n517_), .A3(new_n472_), .A4(new_n382_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n518_), .A3(KEYINPUT20), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n519_), .A2(new_n442_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n495_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n491_), .A2(new_n500_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n495_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n502_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT27), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT96), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n511_), .B2(new_n472_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(new_n390_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n470_), .A2(new_n530_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n529_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n499_), .B1(new_n534_), .B2(KEYINPUT97), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n447_), .B1(new_n470_), .B2(new_n530_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n512_), .A2(KEYINPUT96), .ZN(new_n537_));
  OAI211_X1 g336(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n441_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n519_), .A2(new_n442_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n495_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT98), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n501_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT98), .B1(new_n520_), .B2(new_n495_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT27), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n528_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT99), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n501_), .A2(new_n544_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n520_), .A2(KEYINPUT98), .A3(new_n495_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n527_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT20), .B1(new_n536_), .B2(new_n537_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n499_), .A3(new_n538_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n541_), .B1(new_n557_), .B2(new_n441_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n553_), .B1(new_n558_), .B2(new_n495_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(KEYINPUT99), .A3(new_n528_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n437_), .B1(new_n550_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G71gat), .B(G99gat), .ZN(new_n562_));
  INV_X1    g361(.A(G43gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n489_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G127gat), .B(G134gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G113gat), .B(G120gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n565_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G227gat), .A2(G233gat), .ZN(new_n571_));
  INV_X1    g370(.A(G15gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT30), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT31), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n570_), .B(new_n575_), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n401_), .A2(new_n406_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n411_), .A2(new_n413_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n569_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n414_), .A2(new_n568_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(KEYINPUT4), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G225gat), .A2(G233gat), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n568_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT4), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n583_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n577_), .A2(new_n578_), .A3(new_n568_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(new_n584_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n583_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G1gat), .B(G29gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G57gat), .B(G85gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n582_), .A2(new_n586_), .B1(new_n589_), .B2(new_n583_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n576_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n601_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n559_), .A2(new_n437_), .A3(new_n603_), .A4(new_n528_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n526_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT95), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n587_), .A2(new_n590_), .A3(new_n596_), .A4(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n580_), .A2(G225gat), .A3(new_n581_), .A4(G233gat), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n588_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n583_), .B1(new_n580_), .B2(KEYINPUT4), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n609_), .B(new_n597_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n607_), .B1(new_n599_), .B2(new_n596_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n495_), .A2(KEYINPUT32), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n554_), .A2(new_n555_), .B1(new_n489_), .B2(new_n390_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n496_), .B1(new_n617_), .B2(new_n538_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n618_), .B2(new_n541_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n523_), .A2(new_n616_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n605_), .A2(new_n615_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n604_), .B1(new_n622_), .B2(new_n437_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n561_), .A2(new_n602_), .B1(new_n623_), .B2(new_n576_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G169gat), .B(G197gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  NAND2_X1  g426(.A1(new_n277_), .A2(new_n241_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n275_), .A2(new_n209_), .A3(new_n276_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(KEYINPUT81), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT81), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n277_), .A2(new_n631_), .A3(new_n241_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n630_), .A2(G229gat), .A3(G233gat), .A4(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n210_), .A2(new_n277_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(new_n629_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT82), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n627_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n627_), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT82), .B(new_n640_), .C1(new_n633_), .C2(new_n636_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n624_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n371_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  AOI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(KEYINPUT100), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n601_), .A3(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(KEYINPUT100), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n264_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n624_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n328_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n370_), .A2(new_n643_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n269_), .B1(new_n656_), .B2(new_n601_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT101), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n651_), .A2(new_n658_), .ZN(G1324gat));
  INV_X1    g458(.A(new_n560_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT99), .B1(new_n559_), .B2(new_n528_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n646_), .A2(new_n270_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n656_), .A2(new_n662_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n666_));
  AND4_X1   g465(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .A4(G8gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n270_), .B1(KEYINPUT102), .B2(KEYINPUT39), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n665_), .A2(new_n668_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n663_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g470(.A(new_n576_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n572_), .B1(new_n656_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT41), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n646_), .A2(new_n572_), .A3(new_n672_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n656_), .A2(new_n437_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G22gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT42), .ZN(new_n679_));
  INV_X1    g478(.A(new_n437_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n680_), .A2(G22gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n645_), .B2(new_n681_), .ZN(G1327gat));
  NOR2_X1   g481(.A1(new_n654_), .A2(new_n264_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR4_X1   g483(.A1(new_n624_), .A2(new_n684_), .A3(new_n370_), .A4(new_n643_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n686_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n689_), .A2(G29gat), .A3(new_n603_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n680_), .B(new_n602_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n437_), .A2(new_n603_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n548_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n615_), .A2(new_n605_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n619_), .A2(new_n621_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n437_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n576_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n692_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n691_), .B1(new_n699_), .B2(new_n267_), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT43), .B(new_n266_), .C1(new_n692_), .C2(new_n698_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n655_), .A2(new_n328_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n601_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n690_), .B1(new_n707_), .B2(G29gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT104), .ZN(G1328gat));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n687_), .A2(new_n710_), .A3(new_n662_), .A4(new_n688_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT45), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n706_), .A2(new_n662_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n710_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n712_), .B(KEYINPUT46), .C1(new_n713_), .C2(new_n710_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  NAND3_X1  g517(.A1(new_n706_), .A2(G43gat), .A3(new_n672_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n563_), .B1(new_n689_), .B2(new_n576_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n680_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n687_), .A2(new_n437_), .A3(new_n688_), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n706_), .A2(new_n724_), .B1(new_n723_), .B2(new_n725_), .ZN(G1331gat));
  INV_X1    g525(.A(new_n370_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n727_), .A2(new_n328_), .A3(new_n642_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n653_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n603_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n330_), .A2(new_n727_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n624_), .A2(new_n642_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n601_), .A2(new_n294_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1332gat));
  INV_X1    g535(.A(new_n734_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n292_), .A3(new_n662_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n729_), .A2(new_n662_), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT105), .B(KEYINPUT48), .Z(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(G64gat), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n739_), .B2(G64gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT106), .ZN(G1333gat));
  AOI21_X1  g543(.A(new_n283_), .B1(new_n729_), .B2(new_n672_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT49), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n737_), .A2(new_n283_), .A3(new_n672_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n729_), .A2(new_n437_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G78gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n737_), .A2(new_n285_), .A3(new_n437_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT107), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n727_), .A2(new_n684_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n733_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n601_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n328_), .A2(new_n643_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n370_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT108), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n370_), .A2(new_n763_), .A3(new_n760_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT43), .B1(new_n624_), .B2(new_n266_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n699_), .A2(new_n691_), .A3(new_n267_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n762_), .A2(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n601_), .A2(G85gat), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT109), .Z(new_n769_));
  AOI21_X1  g568(.A(new_n758_), .B1(new_n767_), .B2(new_n769_), .ZN(G1336gat));
  INV_X1    g569(.A(new_n662_), .ZN(new_n771_));
  OR3_X1    g570(.A1(new_n756_), .A2(G92gat), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n763_), .B1(new_n370_), .B2(new_n760_), .ZN(new_n773_));
  AOI211_X1 g572(.A(KEYINPUT108), .B(new_n759_), .C1(new_n365_), .C2(new_n369_), .ZN(new_n774_));
  OAI22_X1  g573(.A1(new_n700_), .A2(new_n701_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G92gat), .B1(new_n775_), .B2(new_n771_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n776_), .ZN(G1337gat));
  AND4_X1   g576(.A1(new_n672_), .A2(new_n757_), .A3(new_n220_), .A4(new_n222_), .ZN(new_n778_));
  INV_X1    g577(.A(G99gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n767_), .B2(new_n672_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781_));
  OAI22_X1  g580(.A1(new_n778_), .A2(new_n780_), .B1(new_n781_), .B2(KEYINPUT51), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(KEYINPUT51), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(G1338gat));
  NOR3_X1   g583(.A1(new_n756_), .A2(G106gat), .A3(new_n680_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n762_), .A2(new_n764_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n765_), .A2(new_n766_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .A4(new_n437_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(G106gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT111), .B1(new_n775_), .B2(new_n680_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n787_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(new_n787_), .A3(G106gat), .A4(new_n791_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n786_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT113), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n791_), .A2(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n790_), .B1(new_n767_), .B2(new_n437_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT52), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n795_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n786_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n798_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n805_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n803_), .B1(new_n802_), .B2(new_n786_), .ZN(new_n808_));
  AOI211_X1 g607(.A(KEYINPUT113), .B(new_n785_), .C1(new_n801_), .C2(new_n795_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n810_), .ZN(G1339gat));
  NAND3_X1  g610(.A1(new_n561_), .A2(new_n601_), .A3(new_n672_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n345_), .A2(new_n814_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n815_), .A2(KEYINPUT114), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(KEYINPUT114), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n333_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n346_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n345_), .A2(new_n814_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n816_), .A2(new_n817_), .A3(new_n819_), .A4(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n353_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(KEYINPUT56), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n821_), .A2(KEYINPUT115), .A3(new_n826_), .A4(new_n822_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n825_), .A2(new_n642_), .A3(new_n358_), .A4(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n633_), .A2(new_n636_), .A3(new_n627_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n635_), .B1(new_n634_), .B2(new_n629_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n630_), .A2(new_n632_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n635_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n829_), .B1(new_n832_), .B2(new_n627_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n828_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n264_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n652_), .B1(new_n828_), .B2(new_n835_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT57), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n813_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n813_), .B1(new_n840_), .B2(KEYINPUT57), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n821_), .A2(new_n826_), .A3(new_n822_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n833_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n826_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n267_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n849_), .A2(KEYINPUT117), .A3(new_n267_), .A4(new_n850_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n843_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n328_), .B1(new_n842_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n371_), .A2(new_n643_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT54), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n812_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n642_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n812_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n840_), .B(new_n838_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n654_), .B1(new_n864_), .B2(new_n851_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n866_), .B2(new_n858_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n856_), .A2(new_n858_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n861_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n869_), .B2(KEYINPUT59), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n642_), .A2(G113gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT118), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n860_), .B1(new_n870_), .B2(new_n872_), .ZN(G1340gat));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n857_), .B(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n865_), .ZN(new_n876_));
  OAI22_X1  g675(.A1(new_n859_), .A2(new_n862_), .B1(new_n876_), .B2(new_n863_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G120gat), .B1(new_n877_), .B2(new_n727_), .ZN(new_n878_));
  INV_X1    g677(.A(G120gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n727_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n859_), .B(new_n880_), .C1(KEYINPUT60), .C2(new_n879_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(G1341gat));
  AOI211_X1 g681(.A(new_n328_), .B(new_n812_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT119), .B1(new_n883_), .B2(G127gat), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885_));
  INV_X1    g684(.A(G127gat), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n885_), .B(new_n886_), .C1(new_n869_), .C2(new_n328_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n328_), .A2(new_n886_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n884_), .A2(new_n887_), .B1(new_n870_), .B2(new_n888_), .ZN(G1342gat));
  OAI21_X1  g688(.A(G134gat), .B1(new_n877_), .B2(new_n266_), .ZN(new_n890_));
  OR3_X1    g689(.A1(new_n869_), .A2(G134gat), .A3(new_n264_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1343gat));
  NAND4_X1  g691(.A1(new_n771_), .A2(new_n601_), .A3(new_n437_), .A4(new_n576_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT120), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n868_), .A2(new_n642_), .A3(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g695(.A1(new_n868_), .A2(new_n370_), .A3(new_n894_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT121), .B(G148gat), .ZN(new_n898_));
  XOR2_X1   g697(.A(new_n897_), .B(new_n898_), .Z(G1345gat));
  NAND3_X1  g698(.A1(new_n868_), .A2(new_n654_), .A3(new_n894_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  NAND2_X1  g701(.A1(new_n868_), .A2(new_n894_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G162gat), .B1(new_n903_), .B2(new_n266_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n264_), .A2(G162gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n903_), .B2(new_n905_), .ZN(G1347gat));
  NAND2_X1  g705(.A1(new_n662_), .A2(new_n602_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n876_), .A2(new_n437_), .A3(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT22), .B(G169gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n642_), .A2(new_n909_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT123), .Z(new_n911_));
  NAND2_X1  g710(.A1(new_n908_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n907_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n642_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT122), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n680_), .B(new_n915_), .C1(new_n875_), .C2(new_n865_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(new_n917_), .A3(G169gat), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n916_), .B2(G169gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n912_), .B1(new_n919_), .B2(new_n920_), .ZN(G1348gat));
  NAND2_X1  g720(.A1(new_n908_), .A2(new_n370_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n437_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n727_), .A2(new_n465_), .A3(new_n907_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n922_), .A2(new_n465_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NOR3_X1   g724(.A1(new_n907_), .A2(new_n448_), .A3(new_n328_), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n680_), .B(new_n926_), .C1(new_n875_), .C2(new_n865_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT124), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n907_), .A2(new_n328_), .ZN(new_n929_));
  AOI21_X1  g728(.A(G183gat), .B1(new_n923_), .B2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n908_), .A2(new_n449_), .A3(new_n652_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n908_), .A2(new_n267_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n460_), .ZN(G1351gat));
  NAND4_X1  g733(.A1(new_n662_), .A2(new_n603_), .A3(new_n437_), .A4(new_n576_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n642_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n370_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n372_), .A2(KEYINPUT125), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n939_), .B(new_n940_), .ZN(G1353gat));
  OR2_X1    g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  AND4_X1   g742(.A1(new_n654_), .A2(new_n936_), .A3(new_n942_), .A4(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n942_), .B1(new_n936_), .B2(new_n654_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1354gat));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT126), .B(G218gat), .Z(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n936_), .B2(new_n652_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n267_), .A2(new_n948_), .ZN(new_n950_));
  AOI211_X1 g749(.A(new_n935_), .B(new_n950_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n947_), .B1(new_n949_), .B2(new_n951_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n936_), .A2(new_n267_), .A3(new_n948_), .ZN(new_n953_));
  AOI211_X1 g752(.A(new_n264_), .B(new_n935_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n954_));
  OAI211_X1 g753(.A(new_n953_), .B(KEYINPUT127), .C1(new_n954_), .C2(new_n948_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n952_), .A2(new_n955_), .ZN(G1355gat));
endmodule


