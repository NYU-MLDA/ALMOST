//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_;
  INV_X1    g000(.A(KEYINPUT10), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT10), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT64), .B1(new_n203_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(KEYINPUT10), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n215_));
  OR2_X1    g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(KEYINPUT9), .A3(new_n214_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT6), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT6), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n213_), .A2(new_n215_), .A3(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G71gat), .B(G78gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT11), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n226_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n235_));
  OR3_X1    g034(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n222_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238_));
  INV_X1    g037(.A(new_n214_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n216_), .A2(KEYINPUT65), .A3(new_n214_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n237_), .A2(KEYINPUT8), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT8), .ZN(new_n245_));
  INV_X1    g044(.A(new_n243_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n222_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n225_), .B(new_n234_), .C1(new_n244_), .C2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT66), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n225_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n233_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G230gat), .A2(G233gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT8), .B1(new_n237_), .B2(new_n243_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n246_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n223_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n256_), .A2(new_n257_), .B1(new_n258_), .B2(new_n215_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n255_), .B1(new_n259_), .B2(new_n234_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n259_), .B2(new_n234_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n251_), .A2(KEYINPUT12), .A3(new_n233_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n253_), .A2(new_n255_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G120gat), .B(G148gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n265_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT13), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n272_), .A2(new_n273_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G29gat), .B(G36gat), .ZN(new_n277_));
  INV_X1    g076(.A(G43gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G50gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT15), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G50gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n279_), .B(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n284_), .A2(KEYINPUT15), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n251_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G232gat), .A2(G233gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT70), .Z(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT69), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT34), .Z(new_n290_));
  OAI221_X1 g089(.A(new_n286_), .B1(KEYINPUT35), .B2(new_n290_), .C1(new_n251_), .C2(new_n280_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(KEYINPUT35), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n292_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G190gat), .B(G218gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G134gat), .ZN(new_n297_));
  INV_X1    g096(.A(G162gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT36), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n295_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n299_), .B(KEYINPUT36), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n293_), .A2(new_n304_), .A3(new_n294_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT37), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G127gat), .B(G155gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT16), .ZN(new_n309_));
  INV_X1    g108(.A(G183gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G211gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT71), .A3(KEYINPUT17), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G15gat), .B(G22gat), .ZN(new_n315_));
  INV_X1    g114(.A(G1gat), .ZN(new_n316_));
  INV_X1    g115(.A(G8gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT14), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G8gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G231gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(new_n234_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n314_), .A2(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n314_), .B(new_n324_), .C1(KEYINPUT17), .C2(new_n313_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT37), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n302_), .A2(new_n329_), .A3(new_n305_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n307_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G141gat), .ZN(new_n333_));
  INV_X1    g132(.A(G169gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n335_), .B(G197gat), .Z(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n321_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G229gat), .A2(G233gat), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n280_), .A2(new_n321_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT72), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n338_), .A2(new_n343_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n280_), .A2(new_n321_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n339_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n337_), .B1(new_n345_), .B2(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n342_), .A2(new_n349_), .A3(new_n344_), .A4(new_n337_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT73), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(G183gat), .A3(G190gat), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n356_), .A2(KEYINPUT76), .ZN(new_n357_));
  INV_X1    g156(.A(G190gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT23), .B1(new_n310_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(KEYINPUT76), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  OR3_X1    g160(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT75), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n361_), .A2(KEYINPUT77), .A3(new_n362_), .ZN(new_n371_));
  OR3_X1    g170(.A1(new_n310_), .A2(KEYINPUT74), .A3(KEYINPUT25), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT26), .B(G190gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT25), .B1(new_n310_), .B2(KEYINPUT74), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n365_), .A2(new_n370_), .A3(new_n371_), .A4(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n359_), .A2(new_n356_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(G183gat), .B2(G190gat), .ZN(new_n378_));
  INV_X1    g177(.A(G176gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n334_), .B2(KEYINPUT22), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT22), .B(G169gat), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n379_), .B(new_n381_), .C1(new_n382_), .C2(new_n380_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n378_), .A2(new_n367_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n376_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(new_n278_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G71gat), .B(G99gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT30), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G227gat), .A2(G233gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n389_), .B(G15gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n388_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n386_), .B(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n392_), .A2(KEYINPUT80), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(KEYINPUT80), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G127gat), .B(G134gat), .ZN(new_n395_));
  INV_X1    g194(.A(G113gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(G120gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OR3_X1    g201(.A1(new_n393_), .A2(new_n394_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT94), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405_));
  INV_X1    g204(.A(G141gat), .ZN(new_n406_));
  INV_X1    g205(.A(G148gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT2), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G141gat), .A2(G148gat), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n408_), .A2(KEYINPUT3), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT2), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n411_), .B(new_n413_), .C1(KEYINPUT3), .C2(new_n408_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G155gat), .B(G162gat), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G155gat), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n417_), .A2(new_n298_), .A3(KEYINPUT1), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT1), .B1(new_n417_), .B2(new_n298_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n418_), .B(new_n419_), .C1(G155gat), .C2(G162gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G141gat), .A2(G148gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n410_), .A3(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n399_), .A2(new_n404_), .A3(new_n416_), .A4(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n397_), .B(G120gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n416_), .A2(new_n423_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n425_), .B1(new_n426_), .B2(KEYINPUT94), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n424_), .A2(new_n427_), .A3(KEYINPUT4), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT95), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n425_), .A2(new_n426_), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n428_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n424_), .A2(new_n427_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n429_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(KEYINPUT97), .B(G1gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G57gat), .B(G85gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G29gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n440_), .B(new_n442_), .Z(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n434_), .B(new_n443_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n394_), .A2(new_n402_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n403_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n426_), .A2(KEYINPUT29), .ZN(new_n453_));
  XOR2_X1   g252(.A(KEYINPUT84), .B(KEYINPUT21), .Z(new_n454_));
  XNOR2_X1  g253(.A(G197gat), .B(G204gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G211gat), .B(G218gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT21), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(new_n461_), .B2(new_n455_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n458_), .B(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n453_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(G233gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(KEYINPUT83), .A2(G228gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT83), .A2(G228gat), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n465_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n452_), .B1(new_n464_), .B2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n458_), .B(new_n462_), .Z(new_n471_));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n469_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n463_), .A2(KEYINPUT86), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .A4(new_n453_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n463_), .B(new_n472_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n478_), .A2(new_n452_), .A3(new_n474_), .A4(new_n453_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G78gat), .B(G106gat), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT88), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n477_), .A2(new_n479_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n480_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n426_), .A2(KEYINPUT29), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT82), .B(KEYINPUT28), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G22gat), .B(G50gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n426_), .A2(KEYINPUT29), .ZN(new_n491_));
  INV_X1    g290(.A(new_n488_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n489_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n490_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT88), .A4(new_n481_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n484_), .A2(new_n486_), .A3(new_n497_), .A4(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n496_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n502_), .A2(KEYINPUT89), .A3(new_n498_), .A4(new_n484_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n486_), .A2(new_n482_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n501_), .A2(new_n503_), .B1(new_n504_), .B2(new_n496_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n361_), .B1(G183gat), .B2(G190gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n382_), .A2(new_n379_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n361_), .B(KEYINPUT91), .C1(G183gat), .C2(G190gat), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .A4(new_n367_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT25), .B(G183gat), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n373_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n369_), .A2(new_n366_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n377_), .A4(new_n362_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n511_), .A2(new_n471_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n473_), .A2(new_n475_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n385_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT20), .B(new_n517_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G226gat), .A2(G233gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT90), .Z(new_n522_));
  XOR2_X1   g321(.A(new_n522_), .B(KEYINPUT19), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n519_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n511_), .A2(new_n516_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n463_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n523_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n525_), .A2(new_n527_), .A3(KEYINPUT20), .A4(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G8gat), .B(G36gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT18), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G64gat), .B(G92gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n524_), .A2(new_n536_), .A3(new_n529_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT27), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n520_), .A2(new_n528_), .ZN(new_n541_));
  AND4_X1   g340(.A1(KEYINPUT20), .A2(new_n525_), .A3(new_n523_), .A4(new_n527_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n536_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n543_), .A2(new_n538_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n544_), .B2(KEYINPUT27), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT98), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n505_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n505_), .B2(new_n545_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n451_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n403_), .A2(new_n449_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n543_), .A2(new_n538_), .A3(KEYINPUT27), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n538_), .A2(new_n539_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(KEYINPUT27), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n505_), .A2(new_n553_), .A3(new_n447_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n428_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n435_), .B2(new_n430_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT33), .B1(new_n556_), .B2(new_n443_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n446_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT33), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n446_), .A2(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n558_), .A2(new_n538_), .A3(new_n539_), .A4(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT32), .B(new_n537_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n530_), .B1(new_n563_), .B2(new_n536_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n564_), .A3(new_n447_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n505_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n550_), .B1(new_n554_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n354_), .B1(new_n549_), .B2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(KEYINPUT99), .ZN(new_n570_));
  INV_X1    g369(.A(new_n354_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n501_), .A2(new_n503_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n504_), .A2(new_n496_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT98), .B1(new_n574_), .B2(new_n553_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n505_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n450_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n403_), .A2(new_n449_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(new_n448_), .A3(new_n545_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n505_), .A2(new_n566_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n571_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n276_), .B(new_n332_), .C1(new_n570_), .C2(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n585_), .A2(G1gat), .A3(new_n448_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n586_), .A2(KEYINPUT38), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n306_), .B1(new_n549_), .B2(new_n568_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n276_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n353_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n328_), .A3(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(G1gat), .B1(new_n591_), .B2(new_n448_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n586_), .A2(KEYINPUT38), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n592_), .A3(new_n593_), .ZN(G1324gat));
  INV_X1    g393(.A(KEYINPUT40), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n588_), .A2(new_n328_), .A3(new_n553_), .A4(new_n590_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n597_));
  AND3_X1   g396(.A1(new_n596_), .A2(G8gat), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n596_), .B2(G8gat), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n569_), .A2(KEYINPUT99), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n582_), .A2(new_n583_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n589_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n604_), .A2(new_n317_), .A3(new_n553_), .A4(new_n332_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n600_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n601_), .B1(new_n600_), .B2(new_n605_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n595_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n596_), .A2(G8gat), .ZN(new_n610_));
  INV_X1    g409(.A(new_n597_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n596_), .A2(G8gat), .A3(new_n597_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT101), .B1(new_n609_), .B2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n600_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(KEYINPUT40), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n608_), .A2(new_n617_), .ZN(G1325gat));
  OAI21_X1  g417(.A(G15gat), .B1(new_n591_), .B2(new_n550_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT41), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n585_), .A2(G15gat), .A3(new_n550_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1326gat));
  OR3_X1    g421(.A1(new_n585_), .A2(G22gat), .A3(new_n505_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n591_), .A2(new_n505_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G22gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT103), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n627_), .A3(G22gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n626_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n623_), .B1(new_n631_), .B2(new_n632_), .ZN(G1327gat));
  NAND2_X1  g432(.A1(new_n306_), .A2(new_n327_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT104), .ZN(new_n635_));
  AOI211_X1 g434(.A(new_n589_), .B(new_n635_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n447_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n307_), .A2(new_n330_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n638_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT43), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n549_), .A2(new_n568_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n638_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n327_), .A4(new_n590_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(G29gat), .A3(new_n447_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n642_), .B1(new_n641_), .B2(new_n638_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n638_), .ZN(new_n649_));
  AOI211_X1 g448(.A(KEYINPUT43), .B(new_n649_), .C1(new_n549_), .C2(new_n568_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n327_), .B(new_n590_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n637_), .B1(new_n647_), .B2(new_n653_), .ZN(G1328gat));
  INV_X1    g453(.A(KEYINPUT46), .ZN(new_n655_));
  INV_X1    g454(.A(G36gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n635_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n604_), .A2(new_n656_), .A3(new_n553_), .A4(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT45), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n636_), .A2(KEYINPUT45), .A3(new_n656_), .A4(new_n553_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n545_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n656_), .B1(new_n663_), .B2(new_n645_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n655_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n653_), .A2(new_n553_), .A3(new_n645_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(KEYINPUT46), .A3(new_n660_), .A4(new_n661_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(G1329gat));
  NAND2_X1  g468(.A1(new_n636_), .A2(new_n578_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n278_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n653_), .A2(G43gat), .A3(new_n578_), .A4(new_n645_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n671_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1330gat));
  AOI21_X1  g475(.A(G50gat), .B1(new_n636_), .B2(new_n574_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n645_), .A2(G50gat), .A3(new_n574_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n679_), .B2(new_n653_), .ZN(G1331gat));
  INV_X1    g479(.A(new_n353_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n276_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n641_), .A2(new_n332_), .A3(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT106), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n684_), .A2(KEYINPUT107), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(KEYINPUT107), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n447_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(G57gat), .ZN(new_n688_));
  AND4_X1   g487(.A1(new_n328_), .A2(new_n588_), .A3(new_n589_), .A4(new_n354_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n448_), .A2(new_n688_), .ZN(new_n690_));
  AOI22_X1  g489(.A1(new_n687_), .A2(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(G1332gat));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n689_), .B2(new_n553_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT48), .Z(new_n694_));
  NOR2_X1   g493(.A1(new_n545_), .A2(G64gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT108), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n684_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n694_), .A2(new_n697_), .ZN(G1333gat));
  INV_X1    g497(.A(G71gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n689_), .B2(new_n578_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT49), .Z(new_n701_));
  NAND3_X1  g500(.A1(new_n684_), .A2(new_n699_), .A3(new_n578_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1334gat));
  INV_X1    g502(.A(G78gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n689_), .B2(new_n574_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT50), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n574_), .A2(new_n704_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT109), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n684_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(G1335gat));
  NAND3_X1  g509(.A1(new_n641_), .A2(new_n657_), .A3(new_n682_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n711_), .A2(KEYINPUT110), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(KEYINPUT110), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n447_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n682_), .A2(new_n327_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n447_), .A2(G85gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT111), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n715_), .B1(new_n717_), .B2(new_n719_), .ZN(G1336gat));
  AOI21_X1  g519(.A(G92gat), .B1(new_n714_), .B2(new_n553_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n553_), .A2(G92gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n717_), .B2(new_n722_), .ZN(G1337gat));
  NAND2_X1  g522(.A1(new_n578_), .A2(new_n211_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n204_), .B1(new_n717_), .B2(new_n578_), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT112), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n716_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n578_), .B(new_n728_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G99gat), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n711_), .B(KEYINPUT110), .Z(new_n732_));
  OAI211_X1 g531(.A(new_n730_), .B(new_n731_), .C1(new_n732_), .C2(new_n724_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n727_), .A2(new_n733_), .A3(KEYINPUT51), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT51), .B1(new_n727_), .B2(new_n733_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n644_), .A2(new_n574_), .A3(new_n728_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT114), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n737_), .A2(G106gat), .A3(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n738_), .A2(KEYINPUT114), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n714_), .A2(new_n212_), .A3(new_n574_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n741_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n737_), .A2(G106gat), .A3(new_n739_), .A4(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n742_), .A2(new_n745_), .A3(new_n748_), .A4(new_n743_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  NOR4_X1   g549(.A1(new_n571_), .A2(new_n331_), .A3(new_n589_), .A4(KEYINPUT54), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n331_), .A2(new_n589_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n354_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n306_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n265_), .A2(new_n271_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n262_), .A2(new_n260_), .A3(new_n263_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n262_), .A2(new_n260_), .A3(new_n263_), .A4(KEYINPUT55), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n254_), .B1(new_n264_), .B2(new_n250_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT115), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT66), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n249_), .B(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n262_), .A2(new_n263_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n255_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n761_), .A4(new_n762_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n765_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n270_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n271_), .B1(new_n765_), .B2(new_n771_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT116), .B1(new_n777_), .B2(KEYINPUT56), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(KEYINPUT56), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n758_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n338_), .A2(new_n348_), .A3(new_n340_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n347_), .A2(new_n339_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n336_), .A3(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n351_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n272_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT117), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n272_), .A2(new_n785_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT57), .B(new_n756_), .C1(new_n781_), .C2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n779_), .A2(new_n780_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n758_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n790_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n794_), .B1(new_n797_), .B2(new_n306_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n757_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n777_), .A2(KEYINPUT56), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n773_), .A2(new_n775_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(KEYINPUT118), .A3(new_n780_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n804_), .A3(new_n785_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n802_), .A2(new_n804_), .A3(KEYINPUT58), .A4(new_n785_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n638_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n800_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n787_), .B(new_n789_), .C1(new_n810_), .C2(new_n758_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n811_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n756_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n793_), .A2(new_n798_), .A3(new_n809_), .A4(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n755_), .B1(new_n813_), .B2(new_n327_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n550_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n575_), .A2(new_n576_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n447_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n815_), .A2(KEYINPUT120), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT120), .B1(new_n815_), .B2(new_n818_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n681_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n823_));
  NOR4_X1   g622(.A1(new_n814_), .A2(KEYINPUT59), .A3(new_n550_), .A4(new_n817_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n354_), .A2(new_n396_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n821_), .A2(new_n396_), .B1(new_n825_), .B2(new_n826_), .ZN(G1340gat));
  XNOR2_X1  g626(.A(KEYINPUT121), .B(G120gat), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n276_), .B2(KEYINPUT60), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n829_), .A2(KEYINPUT60), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n830_), .B(new_n831_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n823_), .A2(new_n276_), .A3(new_n824_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n829_), .ZN(G1341gat));
  OAI21_X1  g633(.A(new_n328_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n835_));
  INV_X1    g634(.A(G127gat), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n327_), .A2(new_n836_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n835_), .A2(new_n836_), .B1(new_n825_), .B2(new_n837_), .ZN(G1342gat));
  OAI21_X1  g637(.A(new_n306_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n839_));
  INV_X1    g638(.A(G134gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n649_), .A2(new_n840_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n839_), .A2(new_n840_), .B1(new_n825_), .B2(new_n841_), .ZN(G1343gat));
  NAND2_X1  g641(.A1(new_n574_), .A2(new_n545_), .ZN(new_n843_));
  NOR4_X1   g642(.A1(new_n814_), .A2(new_n448_), .A3(new_n578_), .A4(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n681_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n589_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g647(.A1(new_n844_), .A2(new_n328_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT61), .B(G155gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT122), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n849_), .B(new_n852_), .ZN(G1346gat));
  AOI21_X1  g652(.A(G162gat), .B1(new_n844_), .B2(new_n306_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n649_), .A2(new_n298_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n844_), .B2(new_n855_), .ZN(G1347gat));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n813_), .A2(new_n327_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n755_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n574_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n450_), .A2(new_n545_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n681_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT123), .Z(new_n863_));
  AOI21_X1  g662(.A(new_n334_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n857_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n866_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n863_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n814_), .A2(new_n869_), .A3(new_n574_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT125), .B(new_n865_), .C1(new_n870_), .C2(new_n334_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(new_n868_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n860_), .A2(new_n861_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n382_), .A3(new_n681_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(G1348gat));
  NOR2_X1   g675(.A1(new_n873_), .A2(new_n276_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n379_), .ZN(G1349gat));
  NOR2_X1   g677(.A1(new_n873_), .A2(new_n327_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n513_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n879_), .B2(new_n310_), .ZN(G1350gat));
  OAI21_X1  g680(.A(G190gat), .B1(new_n873_), .B2(new_n649_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n306_), .A2(new_n373_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n873_), .B2(new_n883_), .ZN(G1351gat));
  NOR2_X1   g683(.A1(new_n545_), .A2(new_n447_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n814_), .A2(new_n505_), .A3(new_n578_), .A4(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n681_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n589_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n887_), .A2(new_n328_), .A3(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT126), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n893_), .B(new_n896_), .ZN(G1354gat));
  AOI21_X1  g696(.A(G218gat), .B1(new_n887_), .B2(new_n306_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n814_), .A2(new_n578_), .ZN(new_n899_));
  INV_X1    g698(.A(G218gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n649_), .A2(new_n900_), .ZN(new_n901_));
  AND4_X1   g700(.A1(new_n574_), .A2(new_n899_), .A3(new_n885_), .A4(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT127), .B1(new_n898_), .B2(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n899_), .A2(new_n574_), .A3(new_n306_), .A4(new_n885_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n900_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n887_), .A2(new_n901_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n903_), .A2(new_n908_), .ZN(G1355gat));
endmodule


