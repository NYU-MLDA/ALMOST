//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n202_));
  XOR2_X1   g001(.A(G71gat), .B(G78gat), .Z(new_n203_));
  XOR2_X1   g002(.A(G57gat), .B(G64gat), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G57gat), .B(G64gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT66), .ZN(new_n208_));
  AOI211_X1 g007(.A(new_n202_), .B(new_n203_), .C1(new_n206_), .C2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n203_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(new_n208_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(KEYINPUT11), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n202_), .A3(new_n208_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n209_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT9), .ZN(new_n221_));
  XOR2_X1   g020(.A(G85gat), .B(G92gat), .Z(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(KEYINPUT9), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT10), .B(G99gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(G106gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n225_), .A2(KEYINPUT64), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n224_), .A2(new_n227_), .A3(G106gat), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n218_), .B(new_n223_), .C1(new_n226_), .C2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT7), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n217_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT65), .A3(new_n215_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n230_), .B1(new_n237_), .B2(new_n222_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n222_), .A2(new_n230_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n218_), .B2(new_n232_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n229_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT12), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n214_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n242_), .A2(new_n243_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n214_), .A2(new_n241_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n214_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n214_), .A2(new_n241_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n214_), .A2(new_n241_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G120gat), .B(G148gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(G176gat), .B(G204gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  NAND3_X1  g060(.A1(new_n252_), .A2(new_n256_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n252_), .A2(KEYINPUT69), .A3(new_n256_), .A4(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n252_), .A2(new_n256_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n261_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n266_), .A2(KEYINPUT13), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT13), .B1(new_n266_), .B2(new_n269_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT70), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G29gat), .B(G36gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(G43gat), .B(G50gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G43gat), .B(G50gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(G29gat), .B(G36gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT15), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G15gat), .B(G22gat), .ZN(new_n286_));
  INV_X1    g085(.A(G1gat), .ZN(new_n287_));
  INV_X1    g086(.A(G8gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT14), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G1gat), .B(G8gat), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n291_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n285_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n284_), .A2(new_n293_), .A3(new_n292_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G229gat), .A2(G233gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300_));
  INV_X1    g099(.A(new_n284_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n294_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n302_), .B2(new_n296_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n300_), .A3(new_n296_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n304_), .A2(G229gat), .A3(G233gat), .A4(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G113gat), .B(G141gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT79), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G169gat), .B(G197gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n299_), .A2(new_n306_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n214_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n214_), .A2(new_n317_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n294_), .B(KEYINPUT77), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G127gat), .B(G155gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT16), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G183gat), .B(G211gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT17), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT17), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n322_), .A2(new_n333_), .A3(new_n324_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n277_), .A2(new_n316_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n337_));
  XOR2_X1   g136(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n338_));
  NAND2_X1  g137(.A1(G232gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n337_), .B1(new_n340_), .B2(KEYINPUT35), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n285_), .B2(new_n241_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n229_), .B(new_n284_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(KEYINPUT35), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT72), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n346_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G190gat), .B(G218gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT73), .ZN(new_n352_));
  XOR2_X1   g151(.A(G134gat), .B(G162gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(KEYINPUT36), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n354_), .B(KEYINPUT36), .Z(new_n357_));
  NAND3_X1  g156(.A1(new_n347_), .A2(new_n349_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT88), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT90), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT89), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368_));
  INV_X1    g167(.A(G141gat), .ZN(new_n369_));
  INV_X1    g168(.A(G148gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n365_), .B1(new_n367_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT89), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n366_), .B(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(KEYINPUT90), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n364_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n363_), .B(KEYINPUT1), .Z(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n362_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G141gat), .A2(G148gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n380_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G22gat), .B(G50gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G228gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n364_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n367_), .A2(new_n374_), .A3(new_n365_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT90), .B1(new_n377_), .B2(new_n378_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT29), .ZN(new_n401_));
  OR2_X1    g200(.A1(G197gat), .A2(G204gat), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT92), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G197gat), .A2(G204gat), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(KEYINPUT21), .A4(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G211gat), .B(G218gat), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n402_), .A2(new_n404_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n405_), .B(new_n406_), .C1(new_n407_), .C2(KEYINPUT21), .ZN(new_n408_));
  XOR2_X1   g207(.A(G211gat), .B(G218gat), .Z(new_n409_));
  NAND4_X1  g208(.A1(new_n407_), .A2(new_n409_), .A3(new_n403_), .A4(KEYINPUT21), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n394_), .B1(new_n401_), .B2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n387_), .A2(new_n388_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n408_), .A2(new_n410_), .A3(KEYINPUT93), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT93), .B1(new_n408_), .B2(new_n410_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n394_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n393_), .B1(new_n412_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n394_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n411_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n413_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n401_), .A2(new_n394_), .A3(new_n416_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n393_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n426_));
  AND3_X1   g225(.A1(new_n419_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n419_), .B2(new_n425_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n392_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n419_), .A2(new_n425_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n426_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n419_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n391_), .A3(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G169gat), .A2(G176gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT24), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G169gat), .A2(G176gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT25), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT25), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT26), .B(G190gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n439_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT24), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n438_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT23), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(G183gat), .B2(G190gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(KEYINPUT23), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n448_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT81), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(KEYINPUT23), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n449_), .A2(G183gat), .A3(G190gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(KEYINPUT81), .A3(new_n448_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n446_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(KEYINPUT83), .A2(G176gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(KEYINPUT83), .A2(G176gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT22), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n465_), .B2(G169gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT22), .B(G169gat), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n463_), .B(new_n466_), .C1(new_n467_), .C2(new_n464_), .ZN(new_n468_));
  OAI22_X1  g267(.A1(new_n450_), .A2(new_n452_), .B1(G183gat), .B2(G190gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n436_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n460_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT84), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT84), .ZN(new_n473_));
  INV_X1    g272(.A(new_n439_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n445_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n459_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT81), .B1(new_n458_), .B2(new_n448_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n470_), .B(new_n473_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G99gat), .ZN(new_n482_));
  INV_X1    g281(.A(G43gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485_));
  INV_X1    g284(.A(G15gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n484_), .B(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n481_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n481_), .A2(new_n488_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT31), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n481_), .A2(new_n488_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT31), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n481_), .A2(new_n488_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G134gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G127gat), .ZN(new_n497_));
  INV_X1    g296(.A(G127gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G134gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n499_), .A3(KEYINPUT85), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT85), .B1(new_n497_), .B2(new_n499_), .ZN(new_n502_));
  INV_X1    g301(.A(G120gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G113gat), .ZN(new_n504_));
  INV_X1    g303(.A(G113gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G120gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n510_));
  OAI22_X1  g309(.A1(new_n501_), .A2(new_n502_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n497_), .A2(new_n499_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT85), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n505_), .A2(G120gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n503_), .A2(G113gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT86), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n514_), .A2(new_n517_), .A3(new_n500_), .A4(new_n508_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n511_), .B1(new_n518_), .B2(KEYINPUT87), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(KEYINPUT87), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n491_), .A2(new_n495_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n435_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n500_), .A2(new_n514_), .B1(new_n517_), .B2(new_n508_), .ZN(new_n526_));
  AND4_X1   g325(.A1(new_n500_), .A2(new_n514_), .A3(new_n517_), .A4(new_n508_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n518_), .A2(KEYINPUT87), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n529_), .B(new_n530_), .C1(new_n380_), .C2(new_n386_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n511_), .A2(new_n518_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n398_), .A2(new_n399_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G225gat), .A2(G233gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G1gat), .B(G29gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT0), .ZN(new_n537_));
  INV_X1    g336(.A(G57gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G85gat), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n531_), .A2(KEYINPUT4), .A3(new_n533_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT4), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n400_), .A2(new_n521_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n534_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n535_), .B(new_n540_), .C1(new_n541_), .C2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT99), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n531_), .A2(KEYINPUT4), .A3(new_n533_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n544_), .A3(new_n543_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT99), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n535_), .A4(new_n540_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n535_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n539_), .B(new_n219_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n478_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n473_), .B1(new_n460_), .B2(new_n470_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n416_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G226gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(KEYINPUT96), .B(new_n416_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n463_), .A2(new_n467_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n469_), .A2(new_n566_), .A3(new_n436_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n445_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT25), .B(G183gat), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n569_), .A2(KEYINPUT95), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(KEYINPUT95), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n568_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n474_), .A2(new_n458_), .A3(new_n448_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n567_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(new_n411_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT20), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n561_), .A2(new_n564_), .A3(new_n565_), .A4(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G8gat), .B(G36gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G64gat), .B(G92gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n576_), .B1(new_n574_), .B2(new_n411_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n479_), .B2(new_n416_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n564_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n578_), .A2(new_n583_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n561_), .A2(new_n586_), .A3(new_n565_), .A4(new_n577_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n583_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(new_n564_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n578_), .A2(new_n587_), .A3(KEYINPUT100), .A4(new_n583_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n590_), .A2(KEYINPUT27), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n594_), .A2(KEYINPUT27), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n599_), .A2(KEYINPUT101), .A3(new_n595_), .A4(new_n590_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n602_));
  NAND2_X1  g401(.A1(new_n591_), .A2(new_n593_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n583_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n604_), .B2(new_n594_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT103), .B1(new_n601_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT103), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n608_), .B(new_n605_), .C1(new_n598_), .C2(new_n600_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n525_), .B(new_n556_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n555_), .B1(new_n429_), .B2(new_n434_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n601_), .A2(new_n606_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n592_), .A2(KEYINPUT32), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n578_), .A2(new_n614_), .A3(new_n587_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n591_), .A2(new_n593_), .A3(new_n613_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n555_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n548_), .A2(new_n534_), .A3(new_n543_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n531_), .A2(new_n533_), .A3(new_n544_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n553_), .A2(new_n621_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n546_), .A2(new_n619_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n549_), .A2(KEYINPUT33), .A3(new_n535_), .A4(new_n540_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n623_), .A2(new_n604_), .A3(new_n594_), .A4(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n618_), .B1(new_n625_), .B2(KEYINPUT98), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n604_), .A2(new_n594_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n546_), .A2(new_n619_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n622_), .A2(new_n620_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n624_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n627_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n435_), .B1(new_n626_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n612_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n522_), .A2(new_n523_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n360_), .B1(new_n610_), .B2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n336_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n555_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G1gat), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n277_), .A2(new_n316_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n610_), .A2(new_n636_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n350_), .A2(KEYINPUT75), .A3(new_n355_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n358_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT75), .B1(new_n350_), .B2(new_n355_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT37), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT76), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT76), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n649_), .B(KEYINPUT37), .C1(new_n645_), .C2(new_n646_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n359_), .A2(KEYINPUT37), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n335_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n642_), .A2(new_n643_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n642_), .A2(new_n643_), .A3(KEYINPUT104), .A4(new_n654_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n556_), .A2(G1gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n641_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  AND4_X1   g460(.A1(new_n641_), .A2(new_n657_), .A3(new_n658_), .A4(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n640_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT105), .B(new_n640_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1324gat));
  NOR2_X1   g466(.A1(new_n607_), .A2(new_n609_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n336_), .A2(new_n637_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G8gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT106), .B1(new_n670_), .B2(KEYINPUT39), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT39), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n669_), .A2(new_n672_), .A3(new_n673_), .A4(G8gat), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(KEYINPUT39), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n659_), .A2(new_n288_), .A3(new_n668_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1325gat));
  INV_X1    g479(.A(new_n635_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n638_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G15gat), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT41), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(KEYINPUT41), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n681_), .A2(new_n486_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n684_), .B(new_n685_), .C1(new_n655_), .C2(new_n686_), .ZN(G1326gat));
  INV_X1    g486(.A(G22gat), .ZN(new_n688_));
  INV_X1    g487(.A(new_n435_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n638_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT42), .Z(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n688_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT107), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n655_), .B2(new_n693_), .ZN(G1327gat));
  INV_X1    g493(.A(new_n335_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(new_n359_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n642_), .A2(new_n643_), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G29gat), .B1(new_n697_), .B2(new_n555_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n277_), .A2(new_n316_), .A3(new_n695_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n643_), .B2(new_n653_), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT43), .B(new_n652_), .C1(new_n610_), .C2(new_n636_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n705_), .A2(G29gat), .A3(new_n555_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT44), .B(new_n699_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n698_), .B1(new_n706_), .B2(new_n707_), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n668_), .A3(new_n707_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G36gat), .ZN(new_n710_));
  INV_X1    g509(.A(G36gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n697_), .A2(new_n711_), .A3(new_n668_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n710_), .A2(new_n714_), .A3(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1329gat));
  NAND4_X1  g518(.A1(new_n705_), .A2(G43gat), .A3(new_n681_), .A4(new_n707_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n697_), .A2(new_n681_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n483_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1330gat));
  NOR2_X1   g524(.A1(new_n435_), .A2(G50gat), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT111), .Z(new_n727_));
  NAND2_X1  g526(.A1(new_n697_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n705_), .A2(new_n689_), .A3(new_n707_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n729_), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT110), .B1(new_n729_), .B2(G50gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(G1331gat));
  AOI21_X1  g531(.A(new_n315_), .B1(new_n610_), .B2(new_n636_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT112), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(KEYINPUT112), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n276_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(new_n654_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n555_), .ZN(new_n738_));
  AND4_X1   g537(.A1(new_n637_), .A2(new_n316_), .A3(new_n277_), .A4(new_n695_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(G57gat), .A3(new_n555_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT113), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n739_), .B2(new_n668_), .ZN(new_n744_));
  XOR2_X1   g543(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n737_), .A2(new_n743_), .A3(new_n668_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1333gat));
  INV_X1    g547(.A(G71gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n739_), .B2(new_n681_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT49), .Z(new_n751_));
  NAND2_X1  g550(.A1(new_n681_), .A2(new_n749_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT115), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n737_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n754_), .ZN(G1334gat));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n739_), .B2(new_n689_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT50), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n737_), .A2(new_n756_), .A3(new_n689_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1335gat));
  AND2_X1   g559(.A1(new_n736_), .A2(new_n696_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n219_), .A3(new_n555_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n701_), .A2(new_n702_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n276_), .A2(new_n315_), .A3(new_n695_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n555_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n762_), .B1(new_n767_), .B2(new_n219_), .ZN(G1336gat));
  NAND3_X1  g567(.A1(new_n761_), .A2(new_n220_), .A3(new_n668_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n668_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(new_n220_), .ZN(G1337gat));
  NOR2_X1   g571(.A1(new_n635_), .A2(new_n224_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n736_), .A2(new_n696_), .A3(new_n773_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n681_), .B(new_n764_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(G99gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G99gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g579(.A1(new_n435_), .A2(G106gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n736_), .A2(new_n696_), .A3(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n689_), .B(new_n764_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(G106gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n783_), .B2(G106gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g587(.A(new_n316_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n248_), .A2(KEYINPUT55), .A3(new_n250_), .A4(new_n251_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(KEYINPUT119), .A3(new_n253_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n255_), .B1(new_n254_), .B2(new_n246_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n253_), .A2(KEYINPUT119), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n792_), .A2(KEYINPUT55), .A3(new_n248_), .A4(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n252_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n797_), .B2(new_n268_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n268_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n789_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n304_), .A2(new_n305_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n298_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n313_), .C1(new_n298_), .C2(new_n297_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n312_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n800_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT57), .A3(new_n359_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n797_), .A2(new_n268_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n268_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n805_), .B1(new_n814_), .B2(new_n789_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n809_), .B1(new_n815_), .B2(new_n360_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n804_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n799_), .B2(new_n798_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT58), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n814_), .A2(new_n820_), .A3(new_n817_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n652_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n808_), .B(new_n816_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n653_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(KEYINPUT120), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n335_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n331_), .A2(new_n314_), .A3(new_n312_), .A4(new_n334_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n831_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n652_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n832_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT54), .B1(new_n837_), .B2(new_n653_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n832_), .A2(KEYINPUT118), .A3(new_n833_), .A4(new_n652_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n828_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n668_), .A2(new_n524_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n555_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n826_), .A2(new_n808_), .A3(new_n816_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n846_), .A2(KEYINPUT122), .A3(new_n335_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT122), .B1(new_n846_), .B2(new_n335_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n840_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n843_), .A2(KEYINPUT59), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n845_), .A2(KEYINPUT59), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n505_), .B1(new_n851_), .B2(new_n315_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n845_), .A2(KEYINPUT121), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n841_), .A2(new_n844_), .A3(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n316_), .A2(G113gat), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n853_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT123), .B1(new_n852_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n845_), .A2(KEYINPUT59), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n849_), .A2(new_n850_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n315_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G113gat), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n853_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n858_), .A2(new_n865_), .ZN(G1340gat));
  INV_X1    g665(.A(new_n851_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G120gat), .B1(new_n867_), .B2(new_n276_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n853_), .A2(new_n855_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n277_), .A2(new_n870_), .A3(new_n503_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n870_), .B2(new_n503_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n868_), .A2(new_n873_), .ZN(G1341gat));
  OAI21_X1  g673(.A(G127gat), .B1(new_n867_), .B2(new_n335_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n869_), .A2(new_n498_), .A3(new_n695_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1342gat));
  OAI21_X1  g676(.A(G134gat), .B1(new_n867_), .B2(new_n652_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n869_), .A2(new_n496_), .A3(new_n360_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1343gat));
  NOR4_X1   g679(.A1(new_n668_), .A2(new_n556_), .A3(new_n681_), .A4(new_n435_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n841_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n316_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n369_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n276_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n370_), .ZN(G1345gat));
  NOR2_X1   g685(.A1(new_n882_), .A2(new_n335_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT61), .B(G155gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n882_), .B2(new_n652_), .ZN(new_n890_));
  INV_X1    g689(.A(G162gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n360_), .A2(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n882_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1347gat));
  NAND3_X1  g694(.A1(new_n668_), .A2(new_n556_), .A3(new_n681_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n689_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n849_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(new_n467_), .A3(new_n315_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n315_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n900_), .A2(new_n901_), .A3(G169gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n900_), .B2(G169gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n899_), .B1(new_n902_), .B2(new_n903_), .ZN(G1348gat));
  NAND2_X1  g703(.A1(new_n841_), .A2(new_n435_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n277_), .A2(G176gat), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n905_), .A2(new_n896_), .A3(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n898_), .A2(new_n277_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n463_), .ZN(G1349gat));
  OR3_X1    g708(.A1(new_n905_), .A2(new_n335_), .A3(new_n896_), .ZN(new_n910_));
  INV_X1    g709(.A(G183gat), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n695_), .A2(new_n571_), .A3(new_n570_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n910_), .A2(new_n911_), .B1(new_n898_), .B2(new_n912_), .ZN(G1350gat));
  NAND2_X1  g712(.A1(new_n898_), .A2(new_n653_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G190gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n898_), .A2(new_n360_), .A3(new_n445_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1351gat));
  NAND2_X1  g716(.A1(new_n635_), .A2(new_n611_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT125), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n919_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n841_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n315_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g723(.A1(new_n921_), .A2(new_n276_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1353gat));
  AOI21_X1  g726(.A(new_n335_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n922_), .A2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT127), .ZN(new_n931_));
  XOR2_X1   g730(.A(new_n929_), .B(new_n931_), .Z(G1354gat));
  OR3_X1    g731(.A1(new_n921_), .A2(G218gat), .A3(new_n359_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G218gat), .B1(new_n921_), .B2(new_n652_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1355gat));
endmodule


