//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT22), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(G176gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT79), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n206_), .A2(new_n208_), .A3(new_n219_), .A4(new_n209_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n211_), .A2(new_n212_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n215_), .A2(new_n217_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n205_), .A2(new_n209_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(KEYINPUT24), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n212_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n221_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT21), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(KEYINPUT21), .A3(new_n234_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n221_), .A2(KEYINPUT80), .A3(new_n229_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n232_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT20), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n206_), .A2(new_n208_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT88), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT88), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n206_), .A2(new_n208_), .A3(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n209_), .A3(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n218_), .A2(new_n212_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT89), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n223_), .B(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n222_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n258_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n243_), .B1(new_n257_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n204_), .B1(new_n246_), .B2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n223_), .B(KEYINPUT87), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n222_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n254_), .A2(new_n256_), .B1(new_n266_), .B2(new_n258_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n204_), .B1(new_n267_), .B2(new_n243_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n232_), .A2(new_n244_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(new_n242_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G8gat), .B(G36gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT18), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n264_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n276_), .B1(new_n264_), .B2(new_n272_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n202_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n221_), .A2(KEYINPUT80), .A3(new_n229_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT80), .B1(new_n221_), .B2(new_n229_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n242_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n243_), .A2(new_n262_), .A3(new_n253_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(KEYINPUT20), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n204_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n251_), .A2(new_n255_), .A3(new_n252_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n255_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n262_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n242_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n204_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n289_), .A2(KEYINPUT20), .A3(new_n290_), .A4(new_n245_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n276_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n264_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(KEYINPUT27), .A3(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n279_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n299_));
  AND2_X1   g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(G141gat), .B2(G148gat), .ZN(new_n308_));
  INV_X1    g107(.A(G141gat), .ZN(new_n309_));
  INV_X1    g108(.A(G148gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT3), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n306_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n304_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n305_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n303_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n309_), .A2(new_n310_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n314_), .A2(new_n318_), .A3(new_n315_), .A4(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT1), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n299_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR4_X1   g125(.A1(new_n317_), .A2(new_n322_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G22gat), .B(G50gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G78gat), .B(G106gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n311_), .A2(new_n308_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n316_), .B(new_n338_), .C1(new_n305_), .C2(new_n304_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n302_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n322_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n324_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT84), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n242_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n337_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT29), .B1(new_n317_), .B2(new_n322_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT84), .B1(new_n240_), .B2(new_n241_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n336_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n335_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n349_), .A2(KEYINPUT85), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n345_), .A2(new_n348_), .A3(new_n335_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n349_), .B2(KEYINPUT85), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n333_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n348_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n336_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n334_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n356_), .A2(new_n330_), .A3(new_n351_), .A4(new_n332_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n357_), .A2(KEYINPUT86), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(KEYINPUT86), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n353_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n298_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(G15gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT30), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n270_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G71gat), .B(G99gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G43gat), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n368_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G134gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G127gat), .ZN(new_n373_));
  INV_X1    g172(.A(G127gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G134gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G120gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G113gat), .ZN(new_n378_));
  INV_X1    g177(.A(G113gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G120gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n373_), .A2(new_n375_), .A3(new_n378_), .A4(new_n380_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n382_), .A2(new_n383_), .A3(KEYINPUT81), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT81), .B1(new_n382_), .B2(new_n383_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n386_), .B(KEYINPUT31), .Z(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT82), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n371_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n387_), .B(KEYINPUT82), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n369_), .A2(new_n390_), .A3(new_n370_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT93), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT94), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n395_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI22_X1  g201(.A1(new_n384_), .A2(new_n385_), .B1(new_n317_), .B2(new_n322_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n403_), .B2(KEYINPUT4), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n382_), .A2(new_n383_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n340_), .A2(new_n341_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(new_n406_), .A3(KEYINPUT91), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT91), .ZN(new_n408_));
  OAI221_X1 g207(.A(new_n408_), .B1(new_n317_), .B2(new_n322_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n404_), .B1(new_n410_), .B2(KEYINPUT4), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n402_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n400_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n401_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n398_), .B(new_n399_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n414_), .B(new_n415_), .C1(new_n417_), .C2(new_n404_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n393_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n361_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n419_), .ZN(new_n422_));
  AND4_X1   g221(.A1(new_n422_), .A2(new_n360_), .A3(new_n279_), .A4(new_n296_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT96), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n276_), .A2(KEYINPUT32), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n292_), .B2(new_n426_), .ZN(new_n427_));
  AOI211_X1 g226(.A(KEYINPUT96), .B(new_n425_), .C1(new_n285_), .C2(new_n291_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n289_), .A2(KEYINPUT20), .A3(new_n245_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n430_), .A2(new_n204_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n425_), .B(KEYINPUT95), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n419_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT97), .B1(new_n429_), .B2(new_n434_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n413_), .A2(new_n418_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT97), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n436_), .B(new_n437_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n401_), .B1(new_n403_), .B2(KEYINPUT4), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n417_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n401_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n440_), .A2(new_n415_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n418_), .A2(KEYINPUT33), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n410_), .A2(KEYINPUT4), .ZN(new_n444_));
  INV_X1    g243(.A(new_n404_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n442_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n245_), .A2(KEYINPUT20), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n290_), .B1(new_n450_), .B2(new_n289_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n282_), .A2(KEYINPUT20), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n290_), .B1(new_n288_), .B2(new_n242_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n293_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n295_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT90), .B1(new_n277_), .B2(new_n278_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n435_), .A2(new_n438_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n360_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n423_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n421_), .B1(new_n462_), .B2(new_n392_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465_));
  INV_X1    g264(.A(G1gat), .ZN(new_n466_));
  INV_X1    g265(.A(G8gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT14), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n471_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT77), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT15), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n474_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n471_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n471_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n474_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n478_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G113gat), .B(G141gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G169gat), .B(G197gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  NAND3_X1  g289(.A1(new_n480_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n490_), .B1(new_n480_), .B2(new_n487_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n464_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n493_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(KEYINPUT78), .A3(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n463_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT69), .ZN(new_n499_));
  INV_X1    g298(.A(G85gat), .ZN(new_n500_));
  INV_X1    g299(.A(G92gat), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT9), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G85gat), .B(G92gat), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n504_), .B2(KEYINPUT64), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G106gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT10), .B(G99gat), .Z(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT64), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n503_), .A2(new_n512_), .A3(KEYINPUT9), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n505_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT66), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n508_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n506_), .B(KEYINPUT6), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT66), .ZN(new_n519_));
  INV_X1    g318(.A(G99gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n520_), .B(new_n509_), .C1(new_n521_), .C2(KEYINPUT7), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n523_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n517_), .A2(new_n519_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n515_), .B1(new_n526_), .B2(new_n503_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n518_), .A2(new_n525_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(new_n515_), .A3(new_n503_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n514_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G57gat), .B(G64gat), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n532_), .A2(KEYINPUT11), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(KEYINPUT11), .ZN(new_n534_));
  XOR2_X1   g333(.A(G71gat), .B(G78gat), .Z(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n531_), .A2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(KEYINPUT12), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n518_), .A2(KEYINPUT66), .B1(new_n522_), .B2(new_n524_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n504_), .B1(new_n542_), .B2(new_n517_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n529_), .B1(new_n543_), .B2(new_n515_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(new_n538_), .A3(new_n514_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n540_), .A2(KEYINPUT12), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G230gat), .A2(G233gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n540_), .A2(new_n545_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(new_n548_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G120gat), .B(G148gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G176gat), .B(G204gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n552_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT68), .ZN(new_n560_));
  INV_X1    g359(.A(new_n548_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n541_), .B2(new_n546_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n557_), .B1(new_n562_), .B2(new_n551_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n559_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(KEYINPUT68), .B(new_n557_), .C1(new_n562_), .C2(new_n551_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n564_), .A2(KEYINPUT13), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT13), .B1(new_n564_), .B2(new_n565_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n499_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT34), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n474_), .B(new_n514_), .C1(new_n527_), .C2(new_n530_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n482_), .B1(new_n544_), .B2(new_n514_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT35), .B(new_n570_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n531_), .A2(new_n483_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(KEYINPUT35), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n570_), .A2(KEYINPUT35), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .A4(new_n571_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(KEYINPUT72), .A3(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G190gat), .B(G218gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n574_), .A2(new_n578_), .A3(KEYINPUT72), .A4(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n574_), .A2(new_n578_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT73), .A3(KEYINPUT37), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n587_), .A2(new_n588_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT73), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT75), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n538_), .B(new_n471_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n605_), .A2(new_n606_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n607_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT76), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(KEYINPUT76), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n599_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n564_), .A2(new_n565_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n564_), .A2(KEYINPUT13), .A3(new_n565_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(KEYINPUT69), .A3(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n568_), .A2(new_n619_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n498_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n498_), .A2(KEYINPUT98), .A3(new_n625_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n466_), .A3(new_n419_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n632_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n463_), .A2(new_n596_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n614_), .ZN(new_n636_));
  AND4_X1   g435(.A1(new_n497_), .A2(new_n568_), .A3(new_n624_), .A4(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT99), .Z(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(new_n419_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n633_), .B(new_n634_), .C1(new_n640_), .C2(new_n466_), .ZN(G1324gat));
  NAND4_X1  g440(.A1(new_n637_), .A2(new_n298_), .A3(new_n463_), .A4(new_n596_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G8gat), .B1(new_n642_), .B2(new_n643_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT39), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n642_), .A2(new_n643_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(G8gat), .A4(new_n644_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n297_), .A2(G8gat), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n628_), .A2(new_n629_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT102), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n651_), .A2(new_n657_), .A3(new_n654_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n659_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n657_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT102), .B(new_n653_), .C1(new_n647_), .C2(new_n650_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n660_), .A2(new_n664_), .ZN(G1325gat));
  AOI21_X1  g464(.A(new_n363_), .B1(new_n639_), .B2(new_n392_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT41), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n630_), .A2(new_n363_), .A3(new_n392_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1326gat));
  INV_X1    g468(.A(G22gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n639_), .B2(new_n360_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT42), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n630_), .A2(new_n670_), .A3(new_n360_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1327gat));
  INV_X1    g473(.A(new_n568_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n624_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n618_), .A2(new_n593_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n498_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n419_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n568_), .A2(new_n624_), .A3(new_n497_), .A4(new_n618_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n594_), .A2(new_n598_), .A3(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n594_), .B2(new_n598_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n463_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT43), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n463_), .A2(new_n691_), .A3(new_n599_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n684_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n683_), .B1(new_n693_), .B2(KEYINPUT44), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n463_), .A2(new_n691_), .A3(new_n599_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n691_), .B1(new_n463_), .B2(new_n688_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT104), .B(new_n695_), .C1(new_n698_), .C2(new_n684_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n684_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n700_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n690_), .A2(new_n692_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n704_), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n700_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n694_), .A2(new_n699_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n419_), .A2(G29gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n682_), .B1(new_n706_), .B2(new_n707_), .ZN(G1328gat));
  INV_X1    g507(.A(G36gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n706_), .B2(new_n298_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n680_), .A2(G36gat), .A3(new_n297_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT45), .ZN(new_n713_));
  OR3_X1    g512(.A1(new_n710_), .A2(new_n711_), .A3(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n711_), .B1(new_n710_), .B2(new_n713_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  NAND2_X1  g515(.A1(new_n694_), .A2(new_n699_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n703_), .A2(new_n705_), .ZN(new_n718_));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n393_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n718_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n706_), .A2(KEYINPUT106), .A3(new_n720_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n719_), .B1(new_n680_), .B2(new_n393_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n723_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT47), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n723_), .A2(new_n728_), .A3(new_n724_), .A4(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1330gat));
  INV_X1    g529(.A(G50gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n706_), .B2(new_n360_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(KEYINPUT107), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(KEYINPUT107), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n360_), .A2(new_n731_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT108), .Z(new_n736_));
  OAI22_X1  g535(.A1(new_n733_), .A2(new_n734_), .B1(new_n680_), .B2(new_n736_), .ZN(G1331gat));
  INV_X1    g536(.A(new_n677_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n497_), .A2(new_n618_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n635_), .A3(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n741_), .A2(G57gat), .A3(new_n419_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(KEYINPUT109), .A3(new_n619_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744_));
  INV_X1    g543(.A(new_n619_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n677_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n497_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n463_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n743_), .A2(new_n746_), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G57gat), .B1(new_n750_), .B2(new_n419_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT110), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT110), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n742_), .B1(new_n752_), .B2(new_n753_), .ZN(G1332gat));
  INV_X1    g553(.A(G64gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n750_), .A2(new_n755_), .A3(new_n298_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n741_), .A2(new_n298_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G64gat), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT48), .B(new_n755_), .C1(new_n741_), .C2(new_n298_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1333gat));
  OR3_X1    g560(.A1(new_n749_), .A2(G71gat), .A3(new_n393_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n741_), .A2(new_n392_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G71gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G71gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(G1334gat));
  INV_X1    g566(.A(G78gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n750_), .A2(new_n768_), .A3(new_n360_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n741_), .A2(new_n360_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G78gat), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT50), .B(new_n768_), .C1(new_n741_), .C2(new_n360_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1335gat));
  NAND3_X1  g573(.A1(new_n738_), .A2(new_n679_), .A3(new_n748_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT111), .ZN(new_n776_));
  AOI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n419_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n618_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n677_), .A2(new_n497_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n704_), .A2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT112), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n422_), .A2(new_n500_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n777_), .B1(new_n781_), .B2(new_n782_), .ZN(G1336gat));
  AOI21_X1  g582(.A(G92gat), .B1(new_n776_), .B2(new_n298_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n297_), .A2(new_n501_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n781_), .B2(new_n785_), .ZN(G1337gat));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(KEYINPUT51), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n776_), .A2(new_n392_), .A3(new_n510_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G99gat), .B1(new_n780_), .B2(new_n393_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n787_), .A2(KEYINPUT51), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(G1338gat));
  NAND3_X1  g592(.A1(new_n776_), .A2(new_n509_), .A3(new_n360_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n704_), .A2(new_n360_), .A3(new_n779_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(G106gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n795_), .B2(G106gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g599(.A1(new_n361_), .A2(new_n419_), .A3(new_n392_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n497_), .A2(new_n559_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n549_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT55), .B1(new_n562_), .B2(KEYINPUT116), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n541_), .A2(KEYINPUT117), .A3(new_n561_), .A4(new_n546_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n805_), .A2(new_n806_), .A3(new_n808_), .A4(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n557_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n557_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n802_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n484_), .A2(new_n486_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n816_), .A2(KEYINPUT118), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(KEYINPUT118), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n479_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n490_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n492_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n564_), .A2(new_n821_), .A3(new_n565_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n596_), .B1(new_n815_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(KEYINPUT119), .A3(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n821_), .A2(new_n559_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT58), .B1(new_n831_), .B2(KEYINPUT120), .ZN(new_n832_));
  INV_X1    g631(.A(new_n830_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n814_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n557_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n832_), .A2(new_n839_), .A3(new_n599_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT57), .B(new_n596_), .C1(new_n815_), .C2(new_n822_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n614_), .B1(new_n829_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n739_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n739_), .B(KEYINPUT114), .C1(new_n566_), .C2(new_n567_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  INV_X1    g648(.A(new_n599_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT115), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n850_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT54), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n848_), .A2(new_n855_), .A3(new_n849_), .A4(new_n850_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n852_), .A2(new_n854_), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n801_), .B1(new_n843_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n379_), .A3(new_n497_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n840_), .A2(new_n841_), .A3(new_n825_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n618_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n801_), .A2(KEYINPUT59), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n497_), .B(new_n864_), .C1(new_n858_), .C2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n859_), .B1(new_n867_), .B2(new_n379_), .ZN(G1340gat));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n858_), .B2(new_n865_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G120gat), .B1(new_n869_), .B2(new_n677_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n843_), .A2(new_n857_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n801_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n377_), .B1(new_n677_), .B2(KEYINPUT60), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(KEYINPUT60), .B2(new_n377_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(KEYINPUT121), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n873_), .A2(new_n878_), .A3(new_n875_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n870_), .B1(new_n877_), .B2(new_n879_), .ZN(G1341gat));
  OAI21_X1  g679(.A(new_n374_), .B1(new_n873_), .B2(new_n618_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT122), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n883_), .B(new_n374_), .C1(new_n873_), .C2(new_n618_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n869_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n614_), .A2(new_n374_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n882_), .A2(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1342gat));
  OAI21_X1  g686(.A(new_n372_), .B1(new_n873_), .B2(new_n596_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  OAI211_X1 g689(.A(KEYINPUT123), .B(new_n372_), .C1(new_n873_), .C2(new_n596_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n599_), .A2(G134gat), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(KEYINPUT124), .Z(new_n893_));
  AOI22_X1  g692(.A1(new_n890_), .A2(new_n891_), .B1(new_n885_), .B2(new_n893_), .ZN(G1343gat));
  NOR4_X1   g693(.A1(new_n298_), .A2(new_n461_), .A3(new_n422_), .A4(new_n392_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n871_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n747_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n309_), .ZN(G1344gat));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n677_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n310_), .ZN(G1345gat));
  AND2_X1   g699(.A1(new_n871_), .A2(new_n895_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n778_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  AOI21_X1  g703(.A(G162gat), .B1(new_n901_), .B2(new_n593_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n688_), .A2(G162gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n901_), .B2(new_n906_), .ZN(G1347gat));
  NAND3_X1  g706(.A1(new_n420_), .A2(new_n461_), .A3(new_n298_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n857_), .B2(new_n861_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n497_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT126), .Z(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  AOI211_X1 g712(.A(new_n747_), .B(new_n908_), .C1(new_n857_), .C2(new_n861_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n205_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n909_), .B2(new_n497_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n913_), .B1(new_n916_), .B2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n908_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n862_), .A2(new_n915_), .A3(new_n497_), .A4(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(G169gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n922_), .A2(new_n917_), .A3(KEYINPUT62), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n912_), .B1(new_n919_), .B2(new_n923_), .ZN(G1348gat));
  AOI21_X1  g723(.A(G176gat), .B1(new_n909_), .B2(new_n738_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n908_), .B1(new_n843_), .B2(new_n857_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n677_), .A2(new_n209_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(G1349gat));
  INV_X1    g727(.A(new_n909_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n929_), .A2(new_n265_), .A3(new_n614_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G183gat), .B1(new_n926_), .B2(new_n778_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n929_), .B2(new_n850_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n909_), .A2(new_n222_), .A3(new_n593_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1351gat));
  NAND4_X1  g734(.A1(new_n298_), .A2(new_n422_), .A3(new_n360_), .A4(new_n393_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n936_), .B1(new_n843_), .B2(new_n857_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n497_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n738_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(KEYINPUT127), .B(G204gat), .ZN(new_n941_));
  XOR2_X1   g740(.A(new_n940_), .B(new_n941_), .Z(G1353gat));
  OR2_X1    g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  NAND2_X1  g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND4_X1   g743(.A1(new_n636_), .A2(new_n937_), .A3(new_n943_), .A4(new_n944_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n943_), .B1(new_n937_), .B2(new_n636_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1354gat));
  INV_X1    g746(.A(G218gat), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n937_), .A2(new_n948_), .A3(new_n593_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n937_), .A2(new_n599_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n948_), .ZN(G1355gat));
endmodule


