//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n859_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(new_n203_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT83), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT84), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(KEYINPUT84), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT31), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT30), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n216_), .A2(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n219_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT80), .B(KEYINPUT23), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n229_), .A2(new_n230_), .B1(new_n231_), .B2(new_n225_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n224_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n222_), .ZN(new_n237_));
  OAI22_X1  g036(.A1(new_n229_), .A2(new_n230_), .B1(new_n231_), .B2(new_n225_), .ZN(new_n238_));
  OR2_X1    g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n215_), .B1(new_n233_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n229_), .A2(new_n230_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n231_), .A2(new_n225_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(new_n223_), .A3(new_n220_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n238_), .A2(new_n239_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n245_), .B(KEYINPUT30), .C1(new_n246_), .C2(new_n237_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G71gat), .B(G99gat), .ZN(new_n248_));
  INV_X1    g047(.A(G43gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G227gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(G15gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n250_), .B(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n241_), .A2(new_n247_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT82), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n241_), .A2(new_n247_), .A3(new_n256_), .A4(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n241_), .B2(new_n247_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT85), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT85), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(new_n263_), .A3(new_n260_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n214_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n266_));
  AOI211_X1 g065(.A(KEYINPUT85), .B(new_n259_), .C1(new_n255_), .C2(new_n257_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n213_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT86), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G228gat), .A2(G233gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(G211gat), .B(G218gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT89), .B(G197gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(G204gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT90), .ZN(new_n274_));
  INV_X1    g073(.A(G204gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(G197gat), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n274_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n278_));
  OAI211_X1 g077(.A(KEYINPUT21), .B(new_n271_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n272_), .A2(new_n275_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT21), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(G197gat), .B2(G204gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n271_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n273_), .A2(new_n281_), .A3(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT3), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT2), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  OR3_X1    g094(.A1(new_n292_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(G155gat), .B2(G162gat), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT87), .B1(new_n298_), .B2(new_n292_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n292_), .A2(KEYINPUT1), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n289_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(new_n287_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT88), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT88), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n306_), .A3(new_n303_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n295_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n270_), .B(new_n286_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n311_));
  OAI21_X1  g110(.A(new_n286_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n270_), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n310_), .A2(KEYINPUT91), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n307_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n306_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT29), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n270_), .A4(new_n286_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G78gat), .B(G106gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n314_), .A2(new_n321_), .A3(new_n325_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n318_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G22gat), .B(G50gat), .Z(new_n330_));
  OR3_X1    g129(.A1(new_n327_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n330_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n324_), .B(new_n326_), .C1(KEYINPUT93), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n326_), .A2(KEYINPUT93), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n331_), .A2(new_n332_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n326_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n325_), .B1(new_n314_), .B2(new_n321_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n335_), .B(new_n336_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n262_), .A2(new_n264_), .A3(new_n214_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n213_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT86), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n269_), .A2(new_n334_), .A3(new_n339_), .A4(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(new_n334_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n265_), .A2(new_n268_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n207_), .A2(new_n204_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT98), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT98), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n207_), .A2(new_n351_), .A3(new_n204_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(new_n315_), .C1(new_n317_), .C2(new_n316_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n308_), .B2(new_n212_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n318_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n354_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n212_), .A2(new_n358_), .A3(new_n318_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n356_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n357_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G1gat), .B(G29gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(G57gat), .B(G85gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n357_), .B(new_n369_), .C1(new_n360_), .C2(new_n363_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT102), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT102), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n375_), .A3(new_n372_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT19), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n222_), .A2(KEYINPUT94), .A3(KEYINPUT24), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT94), .B1(new_n222_), .B2(KEYINPUT24), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n221_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n238_), .A2(new_n220_), .A3(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT95), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n244_), .A2(new_n239_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT96), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n237_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n244_), .A2(KEYINPUT96), .A3(new_n239_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n385_), .A2(new_n391_), .B1(new_n285_), .B2(new_n279_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n245_), .B1(new_n246_), .B2(new_n237_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT20), .B1(new_n286_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n380_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n385_), .A2(new_n391_), .A3(new_n285_), .A4(new_n279_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n380_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n286_), .A2(new_n393_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n396_), .A2(KEYINPUT20), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT18), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT97), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n395_), .A2(new_n399_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n395_), .B2(new_n399_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n378_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT103), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT103), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n409_), .B(new_n378_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n405_), .A2(new_n378_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n392_), .A2(new_n394_), .A3(new_n380_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n391_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n279_), .A2(new_n285_), .A3(new_n384_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT100), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(KEYINPUT100), .B(KEYINPUT20), .C1(new_n414_), .C2(new_n415_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n398_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n413_), .B1(new_n420_), .B2(new_n380_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n412_), .B1(new_n421_), .B2(new_n404_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n377_), .A2(new_n411_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n348_), .A2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n345_), .A2(new_n269_), .A3(new_n343_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n420_), .A2(new_n380_), .ZN(new_n428_));
  OAI211_X1 g227(.A(KEYINPUT101), .B(new_n427_), .C1(new_n428_), .C2(new_n413_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT101), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n395_), .A2(new_n399_), .A3(new_n426_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n429_), .A2(new_n373_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n372_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n405_), .A2(new_n406_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n372_), .A2(new_n434_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n369_), .B1(new_n355_), .B2(new_n362_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n361_), .A2(new_n356_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n360_), .B2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .A4(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n433_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n425_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n424_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  NAND2_X1  g246(.A1(G99gat), .A2(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT65), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT65), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n451_), .A3(KEYINPUT6), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n450_), .B1(G99gat), .B2(G106gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n448_), .A2(KEYINPUT65), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n447_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G85gat), .B(G92gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT68), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT67), .B(KEYINPUT8), .Z(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n449_), .A2(new_n451_), .A3(KEYINPUT6), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT6), .B1(new_n449_), .B2(new_n451_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT69), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n456_), .A2(new_n465_), .A3(new_n452_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n466_), .A3(new_n447_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT70), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n459_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT8), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n467_), .B2(new_n459_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n461_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G71gat), .B(G78gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(G57gat), .B(G64gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(KEYINPUT11), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT71), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT9), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G85gat), .A3(G92gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT10), .B(G99gat), .ZN(new_n481_));
  OAI221_X1 g280(.A(new_n480_), .B1(new_n458_), .B2(new_n479_), .C1(G106gat), .C2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n456_), .A2(new_n452_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n472_), .A2(new_n478_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n472_), .A2(new_n485_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n478_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n472_), .A2(KEYINPUT72), .A3(new_n478_), .A4(new_n485_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G230gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT64), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n467_), .A2(new_n459_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT70), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(KEYINPUT8), .A3(new_n469_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n484_), .B1(new_n499_), .B2(new_n461_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n495_), .B1(new_n500_), .B2(new_n478_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n503_));
  AOI211_X1 g302(.A(KEYINPUT12), .B(new_n478_), .C1(new_n472_), .C2(new_n485_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n501_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G120gat), .B(G148gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(G176gat), .B(G204gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  NAND3_X1  g309(.A1(new_n496_), .A2(new_n505_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT74), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n496_), .B2(new_n505_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AOI211_X1 g313(.A(KEYINPUT74), .B(new_n510_), .C1(new_n496_), .C2(new_n505_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT75), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT13), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520_));
  INV_X1    g319(.A(G1gat), .ZN(new_n521_));
  INV_X1    g320(.A(G8gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G43gat), .B(G50gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(G29gat), .B(G36gat), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n526_), .B(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n526_), .A2(new_n531_), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n531_), .B(KEYINPUT15), .Z(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n534_), .B2(new_n526_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536_));
  MUX2_X1   g335(.A(new_n532_), .B(new_n535_), .S(new_n536_), .Z(new_n537_));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G169gat), .B(G197gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n537_), .B(new_n540_), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n517_), .A2(new_n518_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n543_), .B(new_n544_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n444_), .A2(new_n519_), .A3(new_n542_), .A4(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n526_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n478_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G127gat), .B(G155gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT16), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT78), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G183gat), .B(G211gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n550_), .B1(new_n551_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(KEYINPUT17), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n550_), .B2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT79), .Z(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT34), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n489_), .A2(new_n534_), .B1(new_n565_), .B2(new_n564_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n472_), .A2(new_n485_), .A3(new_n529_), .A4(new_n530_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n489_), .A2(new_n534_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n564_), .A2(new_n565_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT77), .B1(new_n573_), .B2(new_n566_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT77), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n568_), .A2(new_n575_), .A3(new_n567_), .A4(new_n569_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n570_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G190gat), .B(G218gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT36), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT76), .ZN(new_n586_));
  AOI211_X1 g385(.A(new_n586_), .B(new_n570_), .C1(new_n574_), .C2(new_n576_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n561_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n577_), .A2(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n590_), .B(KEYINPUT37), .C1(new_n577_), .C2(new_n582_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n546_), .A2(new_n560_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n377_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n521_), .A3(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT38), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n519_), .A2(new_n545_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n583_), .A2(new_n587_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n560_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n598_), .A2(new_n600_), .A3(new_n542_), .A4(new_n444_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n377_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n596_), .A2(new_n602_), .ZN(G1324gat));
  NAND2_X1  g402(.A1(new_n411_), .A2(new_n422_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n593_), .A2(new_n522_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G8gat), .B1(new_n601_), .B2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT39), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(KEYINPUT39), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT40), .Z(G1325gat));
  AND2_X1   g410(.A1(new_n269_), .A2(new_n343_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G15gat), .B1(new_n601_), .B2(new_n612_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n613_), .A2(KEYINPUT41), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(KEYINPUT41), .ZN(new_n615_));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n612_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n593_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n615_), .A3(new_n618_), .ZN(G1326gat));
  OAI21_X1  g418(.A(G22gat), .B1(new_n601_), .B2(new_n345_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  INV_X1    g420(.A(G22gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n345_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n593_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(G1327gat));
  NAND2_X1  g424(.A1(new_n599_), .A2(new_n560_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n546_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n594_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n560_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n597_), .A2(new_n629_), .A3(new_n541_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n588_), .A2(new_n591_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n348_), .A2(new_n423_), .B1(new_n425_), .B2(new_n442_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n631_), .B(KEYINPUT43), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n444_), .A2(new_n635_), .A3(new_n592_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n444_), .A2(new_n592_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n631_), .B1(new_n638_), .B2(KEYINPUT43), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n630_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n642_), .A2(G29gat), .A3(new_n594_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n424_), .A2(new_n443_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT104), .B1(new_n644_), .B2(new_n635_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(KEYINPUT44), .A3(new_n630_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n628_), .B1(new_n643_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(G1328gat));
  INV_X1    g449(.A(G36gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n627_), .A2(new_n651_), .A3(new_n604_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT45), .Z(new_n653_));
  NOR2_X1   g452(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n642_), .A2(new_n604_), .A3(new_n647_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G36gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT107), .B1(KEYINPUT106), .B2(KEYINPUT46), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n655_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1329gat));
  INV_X1    g460(.A(new_n627_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n249_), .B1(new_n662_), .B2(new_n612_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n642_), .A2(new_n647_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n346_), .A2(G43gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g466(.A1(new_n662_), .A2(G50gat), .A3(new_n345_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n642_), .A2(KEYINPUT108), .A3(new_n647_), .A4(new_n623_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(G50gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n642_), .A2(new_n623_), .A3(new_n647_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT109), .B1(new_n670_), .B2(new_n673_), .ZN(new_n674_));
  AND4_X1   g473(.A1(KEYINPUT109), .A2(new_n673_), .A3(G50gat), .A4(new_n669_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n668_), .B1(new_n674_), .B2(new_n675_), .ZN(G1331gat));
  AOI21_X1  g475(.A(new_n542_), .B1(new_n519_), .B2(new_n545_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n633_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n600_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G57gat), .B1(new_n680_), .B2(new_n377_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n629_), .A3(new_n632_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n377_), .A2(G57gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(G1332gat));
  OR3_X1    g483(.A1(new_n682_), .A2(G64gat), .A3(new_n606_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G64gat), .B1(new_n680_), .B2(new_n606_), .ZN(new_n686_));
  XOR2_X1   g485(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n686_), .A2(new_n687_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(G1333gat));
  OR3_X1    g489(.A1(new_n682_), .A2(G71gat), .A3(new_n612_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n679_), .A2(new_n600_), .A3(new_n617_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G71gat), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(KEYINPUT49), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(KEYINPUT49), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT111), .ZN(G1334gat));
  OAI21_X1  g496(.A(G78gat), .B1(new_n680_), .B2(new_n345_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n699_));
  OR2_X1    g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n699_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n682_), .A2(G78gat), .A3(new_n345_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(G1335gat));
  NOR2_X1   g502(.A1(new_n678_), .A2(new_n629_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n646_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G85gat), .B1(new_n705_), .B2(new_n377_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n677_), .A2(new_n560_), .A3(new_n599_), .A4(new_n444_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT113), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n377_), .A2(G85gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT114), .ZN(G1336gat));
  OAI21_X1  g510(.A(G92gat), .B1(new_n705_), .B2(new_n606_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n606_), .A2(G92gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n708_), .B2(new_n713_), .ZN(G1337gat));
  INV_X1    g513(.A(new_n708_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n481_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n346_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G99gat), .B1(new_n705_), .B2(new_n612_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g519(.A1(new_n708_), .A2(G106gat), .A3(new_n345_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n646_), .A2(new_n704_), .A3(new_n623_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(G106gat), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n722_), .A3(G106gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT53), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT53), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n721_), .B(new_n728_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1339gat));
  NAND2_X1  g529(.A1(new_n606_), .A2(new_n594_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(new_n347_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT57), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n542_), .A2(new_n511_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT115), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n503_), .A2(new_n504_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n488_), .A2(new_n492_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n495_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT55), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n505_), .A2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT55), .B(new_n501_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n510_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n736_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n735_), .B1(new_n745_), .B2(KEYINPUT56), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n488_), .B(new_n492_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n748_));
  AOI22_X1  g547(.A1(new_n748_), .A2(new_n495_), .B1(new_n505_), .B2(new_n740_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n510_), .B1(new_n749_), .B2(new_n742_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n750_), .B2(new_n736_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n537_), .A2(new_n540_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n535_), .A2(G229gat), .A3(G233gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n532_), .A2(new_n536_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(new_n540_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n752_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n746_), .A2(new_n751_), .B1(new_n516_), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n734_), .B1(new_n757_), .B2(new_n599_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n743_), .A2(new_n744_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n760_));
  INV_X1    g559(.A(new_n735_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n751_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n514_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n515_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n756_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n599_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(KEYINPUT57), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n758_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n511_), .A2(new_n756_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n743_), .A2(KEYINPUT56), .A3(new_n744_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT56), .B1(new_n743_), .B2(new_n744_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(KEYINPUT116), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n750_), .A2(new_n777_), .A3(KEYINPUT56), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n772_), .B(new_n773_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n592_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n750_), .B2(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n775_), .A2(KEYINPUT116), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n774_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n772_), .B1(new_n783_), .B2(new_n773_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n780_), .A2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n560_), .B1(new_n769_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n629_), .A2(new_n588_), .A3(new_n591_), .A4(new_n541_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n597_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n788_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n790_), .A2(KEYINPUT54), .A3(new_n519_), .A4(new_n545_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n733_), .B1(new_n786_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G113gat), .B1(new_n794_), .B2(new_n542_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n758_), .B(new_n768_), .C1(new_n784_), .C2(new_n780_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n792_), .B1(new_n797_), .B2(new_n560_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n798_), .B2(new_n733_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT57), .B1(new_n766_), .B2(new_n767_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n734_), .B(new_n599_), .C1(new_n762_), .C2(new_n765_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n784_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(new_n592_), .A3(new_n779_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n629_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT59), .B(new_n732_), .C1(new_n805_), .C2(new_n792_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n799_), .A2(new_n806_), .A3(KEYINPUT118), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT118), .B1(new_n799_), .B2(new_n806_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n542_), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(KEYINPUT119), .B2(G113gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n795_), .B1(new_n809_), .B2(new_n811_), .ZN(G1340gat));
  NAND2_X1  g611(.A1(new_n799_), .A2(new_n806_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT120), .B(G120gat), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT60), .B1(new_n597_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n794_), .A2(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n813_), .A2(new_n597_), .A3(new_n817_), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n818_), .A2(new_n814_), .B1(KEYINPUT60), .B2(new_n817_), .ZN(G1341gat));
  AOI21_X1  g618(.A(G127gat), .B1(new_n794_), .B2(new_n629_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n629_), .A2(G127gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n809_), .B2(new_n821_), .ZN(G1342gat));
  AOI211_X1 g621(.A(KEYINPUT121), .B(G134gat), .C1(new_n794_), .C2(new_n599_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n599_), .B(new_n732_), .C1(new_n805_), .C2(new_n792_), .ZN(new_n825_));
  INV_X1    g624(.A(G134gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT122), .B(G134gat), .Z(new_n829_));
  NOR2_X1   g628(.A1(new_n632_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n809_), .B2(new_n830_), .ZN(G1343gat));
  NOR2_X1   g630(.A1(new_n731_), .A2(new_n344_), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT123), .Z(new_n833_));
  NOR2_X1   g632(.A1(new_n798_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n542_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n597_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n629_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT61), .B(G155gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1346gat));
  INV_X1    g640(.A(G162gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n834_), .A2(new_n842_), .A3(new_n599_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n798_), .A2(new_n632_), .A3(new_n833_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1347gat));
  NAND2_X1  g644(.A1(new_n786_), .A2(new_n793_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n604_), .A2(new_n377_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n847_), .A2(new_n623_), .A3(new_n612_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(G169gat), .B1(new_n849_), .B2(new_n541_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n851_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n849_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n542_), .A3(new_n234_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n853_), .A3(new_n855_), .ZN(G1348gat));
  NOR2_X1   g655(.A1(new_n849_), .A2(new_n598_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n235_), .ZN(G1349gat));
  NOR2_X1   g657(.A1(new_n849_), .A2(new_n560_), .ZN(new_n859_));
  MUX2_X1   g658(.A(G183gat), .B(new_n216_), .S(new_n859_), .Z(G1350gat));
  OAI21_X1  g659(.A(G190gat), .B1(new_n849_), .B2(new_n632_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n599_), .A2(new_n217_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n849_), .B2(new_n862_), .ZN(G1351gat));
  NOR2_X1   g662(.A1(new_n847_), .A2(new_n344_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n798_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n542_), .ZN(new_n867_));
  INV_X1    g666(.A(G197gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(KEYINPUT124), .A3(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n868_), .B2(new_n867_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT124), .B1(new_n867_), .B2(new_n868_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1352gat));
  INV_X1    g671(.A(new_n866_), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n873_), .A2(KEYINPUT125), .A3(new_n275_), .A4(new_n598_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT125), .B(G204gat), .Z(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n866_), .B2(new_n597_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1353gat));
  AOI21_X1  g676(.A(new_n560_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n866_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT126), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n879_), .B(new_n881_), .ZN(G1354gat));
  OR3_X1    g681(.A1(new_n873_), .A2(G218gat), .A3(new_n767_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G218gat), .B1(new_n873_), .B2(new_n632_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1355gat));
endmodule


