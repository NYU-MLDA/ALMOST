//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT90), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT85), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT2), .ZN(new_n208_));
  INV_X1    g007(.A(G141gat), .ZN(new_n209_));
  INV_X1    g008(.A(G148gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT86), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT3), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n211_), .A2(KEYINPUT3), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n205_), .B(new_n206_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n206_), .B(KEYINPUT1), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n205_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n209_), .A2(new_n210_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n207_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT88), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT88), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n217_), .A2(new_n224_), .A3(new_n221_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n203_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(KEYINPUT90), .A3(KEYINPUT29), .A4(new_n225_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G197gat), .B(G204gat), .Z(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT21), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G197gat), .B(G204gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT21), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT92), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT92), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT91), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n230_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G78gat), .B(G106gat), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n243_), .B1(new_n250_), .B2(new_n242_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n247_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n245_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n248_), .B1(new_n254_), .B2(new_n251_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G22gat), .B(G50gat), .Z(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n226_), .A2(new_n227_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n256_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n256_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n259_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n253_), .A2(new_n255_), .A3(new_n262_), .A4(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n265_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n249_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n254_), .A2(new_n248_), .A3(new_n251_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G127gat), .B(G134gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(G113gat), .B(G120gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n223_), .A2(new_n225_), .A3(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n222_), .A2(new_n273_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(KEYINPUT4), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n223_), .A2(new_n277_), .A3(new_n225_), .A4(new_n273_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G225gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT94), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n276_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n274_), .A2(new_n275_), .A3(new_n279_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G1gat), .B(G29gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  NAND3_X1  g086(.A1(new_n281_), .A2(new_n282_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G169gat), .ZN(new_n290_));
  INV_X1    g089(.A(G176gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT24), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(KEYINPUT24), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G190gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT82), .B1(new_n302_), .B2(G183gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT25), .B(G183gat), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n301_), .B(new_n303_), .C1(new_n304_), .C2(KEYINPUT82), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT22), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT83), .B1(new_n307_), .B2(G169gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT22), .B(G169gat), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n291_), .B(new_n308_), .C1(new_n309_), .C2(KEYINPUT83), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n298_), .B2(new_n297_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n298_), .B2(new_n297_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n313_), .A3(new_n294_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n306_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G71gat), .B(G99gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G43gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n315_), .B(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G227gat), .A2(G233gat), .ZN(new_n319_));
  INV_X1    g118(.A(G15gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT30), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT84), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n322_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n273_), .B(KEYINPUT31), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n326_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT84), .B1(new_n330_), .B2(new_n323_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n287_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n289_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT96), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n309_), .A2(new_n291_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n294_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT93), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n313_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n299_), .B1(new_n304_), .B2(new_n301_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n295_), .A3(new_n293_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n242_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT20), .ZN(new_n345_));
  INV_X1    g144(.A(new_n315_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n346_), .B2(new_n241_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT19), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT18), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  NAND2_X1  g154(.A1(new_n242_), .A2(new_n315_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n241_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n350_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(KEYINPUT20), .A4(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n351_), .A2(new_n355_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT27), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n356_), .A2(KEYINPUT20), .A3(new_n357_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n350_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n344_), .A2(new_n347_), .A3(new_n358_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n355_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n336_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n355_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n362_), .A2(new_n350_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n364_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n367_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n370_), .A2(KEYINPUT96), .A3(KEYINPUT27), .A4(new_n360_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n351_), .A2(new_n359_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n367_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n360_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n366_), .A2(new_n371_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  AND4_X1   g175(.A1(new_n266_), .A2(new_n270_), .A3(new_n335_), .A4(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n333_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n270_), .A2(new_n266_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n334_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n288_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n378_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n274_), .A2(new_n275_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n287_), .B1(new_n383_), .B2(new_n280_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n276_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n374_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n288_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n281_), .A2(KEYINPUT33), .A3(new_n282_), .A4(new_n287_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n368_), .A2(new_n369_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n392_));
  MUX2_X1   g191(.A(new_n391_), .B(new_n372_), .S(new_n392_), .Z(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n289_), .B2(new_n334_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n270_), .A2(new_n390_), .A3(new_n394_), .A4(new_n266_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n377_), .B1(new_n382_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G15gat), .B(G22gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G1gat), .A2(G8gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT14), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n399_), .B2(KEYINPUT77), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n399_), .A2(KEYINPUT77), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G1gat), .B(G8gat), .ZN(new_n402_));
  OR3_X1    g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G29gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G43gat), .B(G50gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n405_), .B(new_n408_), .Z(new_n409_));
  NAND2_X1  g208(.A1(G229gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n408_), .B(KEYINPUT15), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n405_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n403_), .A2(new_n404_), .A3(new_n408_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n410_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(G113gat), .B(G141gat), .Z(new_n418_));
  XNOR2_X1  g217(.A(G169gat), .B(G197gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n422_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n412_), .A2(new_n416_), .A3(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT98), .B1(new_n396_), .B2(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n268_), .A2(new_n269_), .A3(new_n267_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n253_), .A2(new_n255_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n381_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n395_), .A3(new_n333_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n377_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT98), .ZN(new_n434_));
  INV_X1    g233(.A(new_n426_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n427_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G230gat), .A2(G233gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(G71gat), .B(G78gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(G57gat), .B(G64gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n439_), .B1(KEYINPUT11), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT68), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT11), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n440_), .B2(KEYINPUT11), .ZN(new_n444_));
  OR3_X1    g243(.A1(new_n441_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n441_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  OAI22_X1  g248(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G99gat), .A2(G106gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(G99gat), .B2(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n450_), .B(new_n453_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G85gat), .ZN(new_n459_));
  INV_X1    g258(.A(G92gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT8), .B1(new_n458_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n456_), .B(KEYINPUT6), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT9), .ZN(new_n466_));
  AND2_X1   g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n461_), .B(new_n466_), .C1(new_n467_), .C2(KEYINPUT65), .ZN(new_n468_));
  OR2_X1    g267(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT64), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT64), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n469_), .A2(new_n471_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT65), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n461_), .A2(new_n476_), .A3(KEYINPUT9), .A4(new_n462_), .ZN(new_n477_));
  AND4_X1   g276(.A1(new_n465_), .A2(new_n468_), .A3(new_n475_), .A4(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n464_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n458_), .A2(KEYINPUT8), .A3(new_n463_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n449_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n455_), .A2(new_n457_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n453_), .A2(new_n450_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n463_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n465_), .A2(new_n468_), .A3(new_n475_), .A4(new_n477_), .ZN(new_n487_));
  AND4_X1   g286(.A1(new_n449_), .A2(new_n486_), .A3(new_n480_), .A4(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n448_), .B1(new_n481_), .B2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n480_), .A3(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT67), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n486_), .A2(new_n449_), .A3(new_n480_), .A4(new_n487_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n447_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n438_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n448_), .A2(KEYINPUT12), .A3(new_n490_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT69), .B1(new_n489_), .B2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n447_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT69), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT12), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n498_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n438_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n495_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G120gat), .B(G148gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT5), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G176gat), .B(G204gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n506_), .A2(KEYINPUT70), .A3(new_n510_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT70), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n502_), .B1(new_n501_), .B2(KEYINPUT12), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n489_), .A2(KEYINPUT69), .A3(new_n499_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n497_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n494_), .B1(new_n516_), .B2(new_n438_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n510_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n513_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n511_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT71), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(KEYINPUT71), .B(new_n511_), .C1(new_n512_), .C2(new_n519_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT13), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n522_), .A2(KEYINPUT13), .A3(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n413_), .A2(new_n490_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(KEYINPUT74), .Z(new_n530_));
  NAND3_X1  g329(.A1(new_n491_), .A2(new_n408_), .A3(new_n492_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n533_));
  NAND2_X1  g332(.A1(G232gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n536_));
  AND2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT76), .B1(new_n535_), .B2(new_n536_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n539_), .A2(new_n529_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n532_), .A2(new_n537_), .B1(new_n531_), .B2(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT36), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT75), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G134gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G162gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n541_), .A2(KEYINPUT36), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT37), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G127gat), .B(G155gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n560_), .B(KEYINPUT17), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n405_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(new_n447_), .ZN(new_n566_));
  MUX2_X1   g365(.A(new_n562_), .B(new_n563_), .S(new_n566_), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT79), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n528_), .A2(new_n555_), .A3(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n437_), .A2(KEYINPUT99), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT99), .B1(new_n437_), .B2(new_n569_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n202_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n396_), .A2(KEYINPUT98), .A3(new_n426_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n434_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n569_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n437_), .A2(KEYINPUT99), .A3(new_n569_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(KEYINPUT100), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n380_), .A2(new_n288_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(G1gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n572_), .A2(new_n579_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT38), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n572_), .A2(new_n579_), .A3(KEYINPUT38), .A4(new_n582_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n528_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n587_), .A2(KEYINPUT101), .A3(new_n435_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT101), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n528_), .B2(new_n426_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n433_), .A2(new_n551_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n567_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n580_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(G1gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n585_), .A2(new_n586_), .A3(new_n596_), .ZN(G1324gat));
  NOR2_X1   g396(.A1(new_n376_), .A2(G8gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n572_), .A2(new_n579_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n376_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n593_), .A2(new_n590_), .A3(new_n600_), .A4(new_n588_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n602_));
  AND3_X1   g401(.A1(new_n601_), .A2(G8gat), .A3(new_n602_), .ZN(new_n603_));
  OR2_X1    g402(.A1(KEYINPUT102), .A2(KEYINPUT39), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n601_), .B2(G8gat), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n599_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n599_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1325gat));
  NAND4_X1  g411(.A1(new_n577_), .A2(new_n320_), .A3(new_n378_), .A4(new_n578_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n594_), .A2(new_n378_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n614_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT41), .B1(new_n614_), .B2(G15gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n613_), .B1(new_n615_), .B2(new_n616_), .ZN(G1326gat));
  INV_X1    g416(.A(G22gat), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n577_), .A2(new_n618_), .A3(new_n379_), .A4(new_n578_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT42), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n594_), .A2(new_n379_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(G22gat), .ZN(new_n622_));
  AOI211_X1 g421(.A(KEYINPUT42), .B(new_n618_), .C1(new_n594_), .C2(new_n379_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n619_), .B1(new_n622_), .B2(new_n623_), .ZN(G1327gat));
  INV_X1    g423(.A(new_n568_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n528_), .A2(new_n625_), .A3(new_n551_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n437_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n581_), .A2(G29gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT105), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n552_), .A2(new_n554_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n625_), .B1(new_n632_), .B2(KEYINPUT43), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n634_), .B1(new_n396_), .B2(new_n631_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n633_), .A2(new_n590_), .A3(new_n588_), .A4(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT44), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n433_), .A2(KEYINPUT43), .A3(new_n555_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n635_), .A2(new_n639_), .A3(new_n568_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n591_), .A3(KEYINPUT44), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n641_), .A3(new_n580_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G29gat), .B1(new_n642_), .B2(new_n643_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n630_), .B1(new_n644_), .B2(new_n645_), .ZN(G1328gat));
  NAND3_X1  g445(.A1(new_n638_), .A2(new_n641_), .A3(new_n600_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G36gat), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n376_), .A2(G36gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n437_), .A2(new_n626_), .A3(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n648_), .A2(KEYINPUT46), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1329gat));
  NAND3_X1  g456(.A1(new_n638_), .A2(new_n641_), .A3(new_n378_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G43gat), .ZN(new_n659_));
  INV_X1    g458(.A(G43gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n627_), .A2(new_n660_), .A3(new_n378_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT47), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n659_), .A2(KEYINPUT47), .A3(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1330gat));
  NAND3_X1  g465(.A1(new_n638_), .A2(new_n641_), .A3(new_n379_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G50gat), .ZN(new_n668_));
  INV_X1    g467(.A(new_n379_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(G50gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT107), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n627_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n668_), .A2(new_n672_), .ZN(G1331gat));
  OAI21_X1  g472(.A(KEYINPUT108), .B1(new_n396_), .B2(new_n435_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n433_), .A2(new_n675_), .A3(new_n426_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n568_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n677_));
  AND4_X1   g476(.A1(new_n528_), .A2(new_n674_), .A3(new_n676_), .A4(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(G57gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n580_), .ZN(new_n680_));
  NOR4_X1   g479(.A1(new_n592_), .A2(new_n587_), .A3(new_n435_), .A4(new_n568_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(new_n580_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n680_), .B1(new_n682_), .B2(new_n679_), .ZN(G1332gat));
  INV_X1    g482(.A(G64gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n681_), .B2(new_n600_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT48), .Z(new_n686_));
  NAND3_X1  g485(.A1(new_n678_), .A2(new_n684_), .A3(new_n600_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1333gat));
  INV_X1    g487(.A(G71gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n681_), .B2(new_n378_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT49), .Z(new_n691_));
  NAND3_X1  g490(.A1(new_n678_), .A2(new_n689_), .A3(new_n378_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1334gat));
  INV_X1    g492(.A(G78gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n681_), .B2(new_n379_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n678_), .A2(new_n694_), .A3(new_n379_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1335gat));
  NOR2_X1   g498(.A1(new_n587_), .A2(new_n435_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n640_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G85gat), .B1(new_n701_), .B2(new_n581_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n551_), .A2(new_n625_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n674_), .A2(new_n676_), .A3(new_n528_), .A4(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n459_), .A3(new_n580_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n702_), .A2(new_n706_), .ZN(G1336gat));
  AOI21_X1  g506(.A(G92gat), .B1(new_n705_), .B2(new_n600_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n701_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n376_), .A2(new_n460_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT110), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n709_), .B2(new_n711_), .ZN(G1337gat));
  NAND4_X1  g511(.A1(new_n705_), .A2(new_n378_), .A3(new_n469_), .A4(new_n474_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n640_), .A2(new_n378_), .A3(new_n700_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(G99gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G99gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT51), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT51), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n720_), .B(new_n713_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1338gat));
  NAND3_X1  g521(.A1(new_n379_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n704_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n640_), .A2(new_n379_), .A3(new_n700_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G106gat), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n726_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n726_), .A2(new_n730_), .A3(new_n731_), .A4(new_n733_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1339gat));
  NOR2_X1   g536(.A1(new_n379_), .A2(new_n600_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n581_), .A2(new_n333_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT57), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n409_), .A2(new_n410_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n414_), .A2(new_n415_), .A3(new_n411_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n422_), .A3(new_n743_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(KEYINPUT119), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n425_), .B1(new_n744_), .B2(KEYINPUT119), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT120), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT116), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n516_), .A2(KEYINPUT116), .A3(new_n438_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n516_), .A2(KEYINPUT55), .A3(new_n438_), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n505_), .B(new_n497_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n756_));
  XOR2_X1   g555(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n754_), .A2(KEYINPUT117), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n516_), .A2(KEYINPUT55), .A3(new_n438_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n757_), .B1(new_n516_), .B2(new_n438_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n504_), .A2(new_n751_), .A3(new_n505_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT116), .B1(new_n516_), .B2(new_n438_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n760_), .B1(new_n763_), .B2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT56), .B(new_n510_), .C1(new_n759_), .C2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT117), .B1(new_n754_), .B2(new_n758_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n763_), .A2(new_n760_), .A3(new_n766_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n518_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n512_), .A2(new_n519_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(new_n426_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n750_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n551_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n741_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n775_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n510_), .B1(new_n759_), .B2(new_n767_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n772_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n779_), .B1(new_n782_), .B2(new_n768_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT57), .B(new_n551_), .C1(new_n783_), .C2(new_n750_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n778_), .A2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n749_), .A2(new_n774_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n769_), .A2(new_n770_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n510_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  AOI211_X1 g588(.A(new_n789_), .B(new_n518_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT58), .B(new_n786_), .C1(new_n788_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n555_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n786_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(KEYINPUT121), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n786_), .C1(new_n788_), .C2(new_n790_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n792_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n567_), .B1(new_n785_), .B2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n677_), .A2(new_n526_), .A3(new_n426_), .A4(new_n527_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n426_), .B(new_n740_), .C1(new_n800_), .C2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT123), .B1(new_n804_), .B2(G113gat), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT123), .ZN(new_n806_));
  INV_X1    g605(.A(G113gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n740_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n806_), .B(new_n807_), .C1(new_n809_), .C2(new_n426_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n568_), .B1(new_n785_), .B2(new_n799_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n803_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n740_), .A2(KEYINPUT59), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n809_), .A2(KEYINPUT59), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n426_), .A2(new_n807_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n805_), .A2(new_n810_), .B1(new_n814_), .B2(new_n815_), .ZN(G1340gat));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n813_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n808_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G120gat), .B1(new_n819_), .B2(new_n587_), .ZN(new_n820_));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n808_), .B(new_n822_), .C1(KEYINPUT60), .C2(new_n821_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1341gat));
  INV_X1    g623(.A(KEYINPUT124), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n568_), .B(new_n740_), .C1(new_n800_), .C2(new_n803_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(G127gat), .ZN(new_n827_));
  INV_X1    g626(.A(G127gat), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT124), .B(new_n828_), .C1(new_n809_), .C2(new_n568_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n567_), .A2(new_n828_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n827_), .A2(new_n829_), .B1(new_n814_), .B2(new_n830_), .ZN(G1342gat));
  OAI21_X1  g630(.A(G134gat), .B1(new_n819_), .B2(new_n631_), .ZN(new_n832_));
  OR3_X1    g631(.A1(new_n809_), .A2(G134gat), .A3(new_n551_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1343gat));
  NAND2_X1  g633(.A1(new_n800_), .A2(new_n803_), .ZN(new_n835_));
  NOR4_X1   g634(.A1(new_n669_), .A2(new_n600_), .A3(new_n581_), .A4(new_n378_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT125), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT125), .ZN(new_n838_));
  INV_X1    g637(.A(new_n836_), .ZN(new_n839_));
  AOI211_X1 g638(.A(new_n838_), .B(new_n839_), .C1(new_n800_), .C2(new_n803_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n435_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G141gat), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n209_), .B(new_n435_), .C1(new_n837_), .C2(new_n840_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1344gat));
  OAI21_X1  g643(.A(new_n528_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(G148gat), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n210_), .B(new_n528_), .C1(new_n837_), .C2(new_n840_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1345gat));
  OAI21_X1  g647(.A(new_n625_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT61), .B(G155gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n850_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n625_), .B(new_n852_), .C1(new_n837_), .C2(new_n840_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1346gat));
  INV_X1    g653(.A(G162gat), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n855_), .B(new_n777_), .C1(new_n837_), .C2(new_n840_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n835_), .A2(new_n836_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n838_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n835_), .A2(KEYINPUT125), .A3(new_n836_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n631_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n856_), .B1(new_n860_), .B2(new_n855_), .ZN(G1347gat));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n600_), .A2(new_n335_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT126), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n379_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n811_), .B2(new_n803_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n435_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n862_), .B1(new_n869_), .B2(new_n290_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n309_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(G1348gat));
  AOI21_X1  g672(.A(G176gat), .B1(new_n867_), .B2(new_n528_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n866_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n587_), .A2(new_n291_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(G1349gat));
  AOI21_X1  g676(.A(G183gat), .B1(new_n875_), .B2(new_n625_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n567_), .A2(new_n304_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n867_), .B2(new_n879_), .ZN(G1350gat));
  NAND3_X1  g679(.A1(new_n867_), .A2(new_n301_), .A3(new_n777_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n867_), .A2(new_n555_), .ZN(new_n882_));
  INV_X1    g681(.A(G190gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1351gat));
  NAND4_X1  g683(.A1(new_n379_), .A2(new_n600_), .A3(new_n581_), .A4(new_n333_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n435_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n528_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g689(.A(new_n567_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT127), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n886_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n893_), .B(new_n894_), .Z(G1354gat));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n886_), .A2(new_n896_), .A3(new_n777_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n886_), .A2(new_n555_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n896_), .ZN(G1355gat));
endmodule


