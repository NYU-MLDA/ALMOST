//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT70), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(new_n204_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(KEYINPUT15), .A3(new_n209_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT72), .B(G15gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(G22gat), .ZN(new_n216_));
  INV_X1    g015(.A(G1gat), .ZN(new_n217_));
  INV_X1    g016(.A(G8gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G1gat), .B(G8gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n221_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n216_), .A2(new_n223_), .A3(new_n219_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n214_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n225_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n210_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n227_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n229_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n225_), .A2(new_n210_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n235_), .A3(KEYINPUT78), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n226_), .A2(new_n230_), .A3(new_n237_), .A4(new_n227_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G113gat), .B(G141gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G169gat), .B(G197gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n240_), .B(new_n241_), .Z(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n236_), .A2(new_n238_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n249_), .B1(G99gat), .B2(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(KEYINPUT6), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n248_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(KEYINPUT6), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(G99gat), .A3(G106gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(KEYINPUT64), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n258_));
  INV_X1    g057(.A(G106gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G85gat), .ZN(new_n262_));
  INV_X1    g061(.A(G92gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G85gat), .A2(G92gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(KEYINPUT9), .A3(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(KEYINPUT9), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n261_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n247_), .B1(new_n257_), .B2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n254_), .A2(new_n255_), .A3(KEYINPUT64), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT64), .B1(new_n254_), .B2(new_n255_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n261_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(KEYINPUT65), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT7), .ZN(new_n277_));
  INV_X1    g076(.A(G99gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n259_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n253_), .A2(new_n282_), .A3(new_n256_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n264_), .A2(new_n265_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n284_), .A2(KEYINPUT8), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n284_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n250_), .A2(new_n252_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n281_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT8), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n276_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n214_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n276_), .A2(new_n229_), .A3(new_n291_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G232gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT34), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT35), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n293_), .A2(new_n294_), .A3(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT69), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n214_), .A2(new_n292_), .B1(new_n298_), .B2(new_n297_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(new_n294_), .ZN(new_n304_));
  OAI22_X1  g103(.A1(new_n301_), .A2(new_n304_), .B1(new_n298_), .B2(new_n297_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(KEYINPUT69), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n297_), .A2(new_n298_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n303_), .A2(new_n302_), .A3(new_n294_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G190gat), .B(G218gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G134gat), .B(G162gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n314_), .A2(KEYINPUT36), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n314_), .A2(KEYINPUT36), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n310_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n317_), .ZN(new_n320_));
  AOI211_X1 g119(.A(KEYINPUT71), .B(new_n320_), .C1(new_n305_), .C2(new_n309_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n316_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT37), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n324_));
  XNOR2_X1  g123(.A(G57gat), .B(G64gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT11), .ZN(new_n326_));
  XOR2_X1   g125(.A(G71gat), .B(G78gat), .Z(new_n327_));
  OR2_X1    g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n325_), .A2(KEYINPUT11), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n327_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n283_), .A2(new_n285_), .B1(new_n289_), .B2(KEYINPUT8), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n332_), .B1(new_n275_), .B2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n291_), .A2(new_n269_), .A3(new_n274_), .A4(new_n331_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT12), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT12), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n337_), .B(new_n332_), .C1(new_n275_), .C2(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G230gat), .A2(G233gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OR4_X1    g140(.A1(KEYINPUT66), .A2(new_n332_), .A3(new_n275_), .A4(new_n333_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n340_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n334_), .A2(KEYINPUT66), .A3(new_n335_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G120gat), .B(G148gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT5), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G176gat), .B(G204gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT67), .B1(new_n347_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n346_), .A2(new_n354_), .A3(new_n351_), .ZN(new_n355_));
  OAI221_X1 g154(.A(new_n324_), .B1(new_n347_), .B2(new_n352_), .C1(new_n353_), .C2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n353_), .A2(new_n355_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n347_), .A2(new_n352_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(KEYINPUT13), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n356_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(G231gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n331_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT73), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(new_n228_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT75), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G127gat), .B(G155gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G183gat), .B(G211gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT17), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n366_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n372_), .A2(new_n373_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n366_), .A2(new_n374_), .A3(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT37), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n316_), .B(new_n381_), .C1(new_n319_), .C2(new_n321_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n323_), .A2(new_n362_), .A3(new_n380_), .A4(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n246_), .B1(new_n383_), .B2(KEYINPUT77), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386_));
  INV_X1    g185(.A(G141gat), .ZN(new_n387_));
  INV_X1    g186(.A(G148gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT2), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G141gat), .A2(G148gat), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n389_), .B(new_n390_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(KEYINPUT85), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT88), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397_));
  OR2_X1    g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT86), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n400_), .A3(KEYINPUT1), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(new_n398_), .C1(KEYINPUT1), .C2(new_n397_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n397_), .B2(KEYINPUT1), .ZN(new_n403_));
  OAI221_X1 g202(.A(new_n394_), .B1(G141gat), .B2(G148gat), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT87), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n399_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G127gat), .B(G134gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G113gat), .B(G120gat), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(KEYINPUT84), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n407_), .A2(new_n408_), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(KEYINPUT4), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n399_), .B(new_n405_), .C1(new_n411_), .C2(new_n409_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(KEYINPUT4), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n416_), .B2(KEYINPUT100), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n413_), .A2(new_n415_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT100), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT4), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n385_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n385_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G85gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT0), .B(G57gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n430_), .A2(KEYINPUT33), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT33), .B(new_n428_), .C1(new_n421_), .C2(new_n423_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT18), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G64gat), .B(G92gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT19), .ZN(new_n440_));
  INV_X1    g239(.A(G183gat), .ZN(new_n441_));
  INV_X1    g240(.A(G190gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT23), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT82), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT23), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(G183gat), .A3(G190gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(G183gat), .B2(G190gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G169gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n443_), .A2(new_n446_), .ZN(new_n451_));
  INV_X1    g250(.A(G169gat), .ZN(new_n452_));
  INV_X1    g251(.A(G176gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n451_), .B1(KEYINPUT24), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT26), .B(G190gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT96), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT25), .B(G183gat), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n455_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT24), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(G169gat), .B2(G176gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n463_), .A2(KEYINPUT97), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n454_), .B(KEYINPUT81), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(KEYINPUT97), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n448_), .A2(new_n450_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G211gat), .B(G218gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT91), .B(G197gat), .ZN(new_n470_));
  INV_X1    g269(.A(G204gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT21), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n473_), .B1(G197gat), .B2(G204gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n469_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G197gat), .A2(G204gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT91), .B(G197gat), .Z(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(G204gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n475_), .B1(KEYINPUT21), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(KEYINPUT21), .A3(new_n469_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI211_X1 g281(.A(new_n438_), .B(new_n440_), .C1(new_n468_), .C2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n481_), .B(KEYINPUT92), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT80), .B(G190gat), .Z(new_n485_));
  OAI21_X1  g284(.A(new_n451_), .B1(new_n485_), .B2(G183gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n450_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n465_), .A2(new_n462_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n447_), .B(new_n488_), .C1(KEYINPUT24), .C2(new_n465_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n485_), .B2(KEYINPUT26), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT79), .B1(new_n441_), .B2(KEYINPUT25), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT79), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n459_), .A2(new_n493_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n491_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n487_), .B1(new_n489_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n484_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n483_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT99), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  OAI221_X1 g299(.A(KEYINPUT20), .B1(new_n482_), .B2(new_n468_), .C1(new_n484_), .C2(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n440_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT98), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n502_), .A2(KEYINPUT98), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n437_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n417_), .A2(new_n420_), .A3(new_n385_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n428_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n505_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n510_), .A2(new_n436_), .A3(new_n503_), .A4(new_n500_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n432_), .A2(new_n506_), .A3(new_n509_), .A4(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n424_), .B(new_n429_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n436_), .A2(KEYINPUT32), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n504_), .A2(new_n515_), .A3(new_n505_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n481_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n468_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT20), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT101), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n497_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n520_), .A2(KEYINPUT101), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n440_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n501_), .A2(new_n440_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n516_), .B1(new_n515_), .B2(new_n526_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n431_), .A2(new_n513_), .B1(new_n514_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n529_));
  INV_X1    g328(.A(G233gat), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n530_), .A2(KEYINPUT90), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(KEYINPUT90), .ZN(new_n532_));
  OAI21_X1  g331(.A(G228gat), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n406_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT29), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n534_), .B1(new_n537_), .B2(new_n518_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n484_), .B(new_n533_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G78gat), .B(G106gat), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n529_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT28), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n535_), .A2(new_n544_), .A3(new_n536_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT28), .B1(new_n406_), .B2(KEYINPUT29), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G22gat), .B(G50gat), .Z(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n549_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n550_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n552_), .B1(new_n553_), .B2(new_n547_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n542_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n540_), .A2(new_n541_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n558_), .A2(new_n554_), .A3(new_n551_), .A4(new_n542_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n551_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n540_), .A2(KEYINPUT95), .A3(new_n541_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT95), .B1(new_n540_), .B2(new_n541_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n506_), .A2(new_n511_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT27), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT102), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT102), .ZN(new_n569_));
  AOI211_X1 g368(.A(new_n569_), .B(KEYINPUT27), .C1(new_n506_), .C2(new_n511_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n436_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n511_), .A2(KEYINPUT27), .ZN(new_n572_));
  OAI22_X1  g371(.A1(new_n568_), .A2(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n424_), .B(new_n428_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n574_), .A2(new_n559_), .A3(new_n557_), .A4(new_n563_), .ZN(new_n575_));
  OAI22_X1  g374(.A1(new_n528_), .A2(new_n565_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n412_), .B(KEYINPUT31), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(KEYINPUT83), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G227gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(G15gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT30), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n496_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n578_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G71gat), .B(G99gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G43gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n584_), .B(new_n586_), .Z(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n564_), .A2(new_n587_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n573_), .A2(new_n589_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n576_), .A2(new_n588_), .B1(new_n574_), .B2(new_n590_), .ZN(new_n591_));
  AOI211_X1 g390(.A(new_n384_), .B(new_n591_), .C1(KEYINPUT77), .C2(new_n383_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n217_), .A3(new_n514_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT38), .ZN(new_n594_));
  INV_X1    g393(.A(new_n362_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n246_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n380_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT104), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n322_), .A2(KEYINPUT103), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n322_), .A2(KEYINPUT103), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n591_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n590_), .A2(new_n574_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n572_), .A2(new_n571_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n566_), .A2(new_n567_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n569_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n566_), .A2(KEYINPUT102), .A3(new_n567_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n606_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n564_), .A2(new_n514_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n504_), .A2(new_n505_), .ZN(new_n612_));
  MUX2_X1   g411(.A(new_n612_), .B(new_n526_), .S(new_n515_), .Z(new_n613_));
  NOR2_X1   g412(.A1(new_n430_), .A2(KEYINPUT33), .ZN(new_n614_));
  OAI22_X1  g413(.A1(new_n574_), .A2(new_n613_), .B1(new_n614_), .B2(new_n512_), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n610_), .A2(new_n611_), .B1(new_n615_), .B2(new_n564_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n605_), .B1(new_n616_), .B2(new_n587_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(KEYINPUT104), .A3(new_n602_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n598_), .B1(new_n604_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n574_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n594_), .A2(new_n621_), .ZN(G1324gat));
  NAND3_X1  g421(.A1(new_n592_), .A2(new_n218_), .A3(new_n573_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n619_), .A2(new_n573_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(G8gat), .ZN(new_n626_));
  AOI211_X1 g425(.A(KEYINPUT39), .B(new_n218_), .C1(new_n619_), .C2(new_n573_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g428(.A1(new_n592_), .A2(new_n580_), .A3(new_n587_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G15gat), .B1(new_n620_), .B2(new_n588_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n632_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(G1326gat));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n592_), .A2(new_n636_), .A3(new_n565_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G22gat), .B1(new_n620_), .B2(new_n564_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(KEYINPUT42), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(KEYINPUT42), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n637_), .B1(new_n639_), .B2(new_n640_), .ZN(G1327gat));
  INV_X1    g440(.A(new_n322_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n380_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n597_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n617_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(G29gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n514_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n323_), .A2(new_n382_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT43), .B1(new_n591_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n617_), .A2(new_n651_), .A3(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n380_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n597_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT44), .B1(new_n653_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n658_), .B(new_n655_), .C1(new_n650_), .C2(new_n652_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n657_), .A2(new_n659_), .A3(new_n574_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n647_), .B1(new_n660_), .B2(new_n646_), .ZN(G1328gat));
  INV_X1    g460(.A(new_n645_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n662_), .A2(G36gat), .A3(new_n610_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT45), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n657_), .A2(new_n659_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n573_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n591_), .A2(KEYINPUT43), .A3(new_n649_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n651_), .B1(new_n617_), .B2(new_n648_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n656_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n658_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n656_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n671_), .A2(new_n665_), .A3(new_n573_), .A4(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G36gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n664_), .B1(new_n667_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n664_), .B(KEYINPUT46), .C1(new_n667_), .C2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1329gat));
  NAND3_X1  g478(.A1(new_n666_), .A2(G43gat), .A3(new_n587_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n662_), .A2(new_n588_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(G43gat), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g482(.A1(new_n662_), .A2(G50gat), .A3(new_n564_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n666_), .A2(new_n685_), .A3(new_n565_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G50gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n666_), .B2(new_n565_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1331gat));
  NOR2_X1   g488(.A1(new_n362_), .A2(new_n246_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n380_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n604_), .B2(new_n618_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G57gat), .B1(new_n693_), .B2(new_n574_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n617_), .A2(new_n690_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n323_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n514_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n694_), .A2(new_n699_), .ZN(G1332gat));
  INV_X1    g499(.A(G64gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n692_), .B2(new_n573_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT48), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(new_n701_), .A3(new_n573_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1333gat));
  INV_X1    g504(.A(G71gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n706_), .A3(new_n587_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G71gat), .B1(new_n693_), .B2(new_n588_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT49), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT49), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(G1334gat));
  INV_X1    g510(.A(G78gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n697_), .A2(new_n712_), .A3(new_n565_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n692_), .A2(new_n565_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(G78gat), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G78gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT108), .Z(G1335gat));
  NAND2_X1  g518(.A1(new_n695_), .A2(new_n643_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n262_), .A3(new_n514_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n690_), .A2(new_n654_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT109), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(new_n514_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n726_), .B2(new_n262_), .ZN(G1336gat));
  NAND3_X1  g526(.A1(new_n721_), .A2(new_n263_), .A3(new_n573_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n725_), .A2(new_n573_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n263_), .ZN(G1337gat));
  AND4_X1   g529(.A1(new_n258_), .A2(new_n721_), .A3(new_n260_), .A4(new_n587_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n278_), .B1(new_n724_), .B2(new_n587_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  AOI211_X1 g535(.A(new_n564_), .B(new_n723_), .C1(new_n650_), .C2(new_n652_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n735_), .B(new_n736_), .C1(new_n737_), .C2(new_n259_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n721_), .A2(new_n259_), .A3(new_n565_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n737_), .B2(new_n259_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n724_), .A2(new_n565_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(KEYINPUT110), .A3(G106gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n743_), .A3(KEYINPUT52), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n740_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n740_), .B2(new_n744_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1339gat));
  INV_X1    g547(.A(G113gat), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT54), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n696_), .A2(new_n750_), .A3(new_n596_), .A4(new_n362_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT54), .B1(new_n383_), .B2(new_n246_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n341_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n343_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT112), .B1(new_n757_), .B2(KEYINPUT55), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n336_), .A2(new_n343_), .A3(new_n338_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  AND4_X1   g559(.A1(KEYINPUT113), .A2(new_n339_), .A3(KEYINPUT55), .A4(new_n340_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT113), .B1(new_n757_), .B2(KEYINPUT55), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT56), .B(new_n351_), .C1(new_n760_), .C2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT115), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n339_), .A2(KEYINPUT55), .A3(new_n340_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n757_), .A2(KEYINPUT113), .A3(KEYINPUT55), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n770_), .A2(new_n756_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(KEYINPUT56), .A4(new_n351_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n351_), .B1(new_n760_), .B2(new_n763_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n765_), .A2(new_n773_), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n226_), .A2(new_n232_), .A3(new_n230_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n227_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n244_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n243_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n357_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n777_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n777_), .A2(KEYINPUT58), .A3(new_n782_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n648_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT116), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n785_), .A2(new_n786_), .A3(new_n789_), .A4(new_n648_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n243_), .B(new_n780_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n246_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n776_), .B2(new_n764_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n793_), .B2(KEYINPUT114), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n795_), .B(new_n792_), .C1(new_n764_), .C2(new_n776_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n642_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT57), .B(new_n642_), .C1(new_n794_), .C2(new_n796_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n788_), .A2(new_n790_), .A3(new_n799_), .A4(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n753_), .B1(new_n801_), .B2(new_n654_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n590_), .A2(new_n514_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n749_), .B1(new_n806_), .B2(new_n596_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT117), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT59), .B1(new_n802_), .B2(new_n804_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n802_), .C2(new_n804_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n753_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n799_), .A2(new_n787_), .A3(new_n800_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n654_), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT59), .B(new_n804_), .C1(new_n814_), .C2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT119), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n813_), .A2(new_n821_), .A3(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n596_), .A2(new_n749_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n808_), .B1(new_n824_), .B2(new_n825_), .ZN(G1340gat));
  XOR2_X1   g625(.A(KEYINPUT120), .B(G120gat), .Z(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n819_), .B2(new_n362_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT121), .B1(new_n827_), .B2(KEYINPUT60), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n595_), .B2(new_n831_), .ZN(new_n832_));
  MUX2_X1   g631(.A(new_n830_), .B(KEYINPUT121), .S(new_n832_), .Z(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n806_), .B2(new_n833_), .ZN(G1341gat));
  AOI21_X1  g633(.A(new_n821_), .B1(new_n813_), .B2(new_n818_), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT119), .B(new_n817_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n380_), .A2(G127gat), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n806_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G127gat), .B1(new_n839_), .B2(new_n380_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT122), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n842_));
  INV_X1    g641(.A(new_n840_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n842_), .B(new_n843_), .C1(new_n823_), .C2(new_n837_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(G1342gat));
  OAI21_X1  g644(.A(G134gat), .B1(new_n823_), .B2(new_n649_), .ZN(new_n846_));
  OR3_X1    g645(.A1(new_n806_), .A2(G134gat), .A3(new_n602_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1343gat));
  NOR3_X1   g647(.A1(new_n564_), .A2(new_n574_), .A3(new_n587_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n803_), .A2(new_n610_), .A3(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n596_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(new_n387_), .ZN(G1344gat));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n362_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n388_), .ZN(G1345gat));
  NOR2_X1   g653(.A1(new_n850_), .A2(new_n654_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT61), .B(G155gat), .Z(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT123), .B(KEYINPUT124), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  OAI21_X1  g658(.A(G162gat), .B1(new_n850_), .B2(new_n649_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n602_), .A2(G162gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n850_), .B2(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT125), .ZN(G1347gat));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n814_), .A2(new_n816_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n514_), .A2(new_n588_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n573_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n565_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n865_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n596_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT22), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n864_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G169gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n452_), .B1(new_n870_), .B2(new_n864_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n872_), .B2(new_n874_), .ZN(G1348gat));
  AOI21_X1  g674(.A(KEYINPUT126), .B1(new_n803_), .B2(new_n564_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n802_), .A2(new_n877_), .A3(new_n565_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n876_), .A2(new_n867_), .A3(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(G176gat), .A3(new_n595_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT127), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n881_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n453_), .B1(new_n869_), .B2(new_n362_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .ZN(G1349gat));
  NOR3_X1   g684(.A1(new_n869_), .A2(new_n459_), .A3(new_n654_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n879_), .A2(new_n380_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n441_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n869_), .B2(new_n649_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n603_), .A2(new_n458_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n869_), .B2(new_n890_), .ZN(G1351gat));
  NOR3_X1   g690(.A1(new_n610_), .A2(new_n575_), .A3(new_n587_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n803_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n246_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g695(.A1(new_n893_), .A2(new_n362_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n471_), .ZN(G1353gat));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n380_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  AND2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n899_), .B2(new_n900_), .ZN(G1354gat));
  OAI21_X1  g702(.A(G218gat), .B1(new_n893_), .B2(new_n649_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n602_), .A2(G218gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n893_), .B2(new_n905_), .ZN(G1355gat));
endmodule


