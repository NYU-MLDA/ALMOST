//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT87), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT86), .B(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n207_), .A2(new_n208_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(KEYINPUT23), .B2(new_n208_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(new_n211_), .B2(new_n206_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT22), .B(G169gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(new_n217_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n216_), .A2(new_n217_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT24), .B1(new_n216_), .B2(new_n217_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT84), .A2(G183gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n228_), .B(KEYINPUT25), .Z(new_n229_));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT26), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(G190gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n229_), .B(new_n232_), .C1(new_n230_), .C2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n224_), .A2(KEYINPUT24), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n227_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n221_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G127gat), .B(G134gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G113gat), .B(G120gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT88), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT88), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT30), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT30), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(new_n246_), .A3(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n237_), .A2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n221_), .A2(new_n245_), .A3(new_n236_), .A4(new_n247_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G15gat), .B(G43gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT31), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n250_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n205_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n204_), .A3(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT21), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT92), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n261_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT91), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT21), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n269_), .A2(new_n261_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(KEYINPUT92), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G228gat), .ZN(new_n273_));
  INV_X1    g072(.A(G233gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT90), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT89), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT1), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n279_), .B(new_n280_), .C1(new_n283_), .C2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n278_), .B(KEYINPUT3), .Z(new_n287_));
  XOR2_X1   g086(.A(new_n280_), .B(KEYINPUT2), .Z(new_n288_));
  OAI211_X1 g087(.A(new_n282_), .B(new_n284_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n277_), .B1(new_n290_), .B2(KEYINPUT29), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n272_), .A2(new_n276_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n276_), .B1(new_n272_), .B2(new_n291_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT93), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n294_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT93), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n292_), .ZN(new_n298_));
  INV_X1    g097(.A(G50gat), .ZN(new_n299_));
  OR3_X1    g098(.A1(new_n290_), .A2(KEYINPUT29), .A3(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT28), .B(G22gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n290_), .B2(KEYINPUT29), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n302_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n295_), .A2(new_n298_), .A3(new_n303_), .A4(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G78gat), .B(G106gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n303_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n309_), .A2(new_n297_), .A3(new_n296_), .A4(new_n292_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n308_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n260_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n260_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n307_), .A2(new_n310_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n308_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n318_), .A3(new_n311_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n237_), .A2(new_n272_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT95), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n225_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT25), .B(G183gat), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n323_), .A2(new_n224_), .B1(new_n233_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n212_), .A2(new_n235_), .A3(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n220_), .B1(new_n223_), .B2(new_n213_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n321_), .B(KEYINPUT20), .C1(new_n272_), .C2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n328_), .A2(new_n272_), .A3(KEYINPUT96), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT96), .B1(new_n328_), .B2(new_n272_), .ZN(new_n335_));
  OAI221_X1 g134(.A(KEYINPUT20), .B1(new_n237_), .B2(new_n272_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n333_), .B1(new_n336_), .B2(new_n332_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G92gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT18), .B(G64gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n333_), .B(new_n343_), .C1(new_n336_), .C2(new_n332_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(KEYINPUT97), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT97), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(new_n346_), .A3(new_n341_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT103), .B(KEYINPUT27), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT4), .B1(new_n244_), .B2(new_n290_), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n290_), .A2(KEYINPUT98), .A3(new_n240_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n244_), .A2(new_n290_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT98), .B1(new_n290_), .B2(new_n240_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n350_), .B1(new_n354_), .B2(KEYINPUT4), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT99), .ZN(new_n357_));
  OR3_X1    g156(.A1(new_n355_), .A2(KEYINPUT100), .A3(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n351_), .A2(new_n356_), .A3(new_n352_), .A4(new_n353_), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n359_), .B(KEYINPUT101), .Z(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT100), .B1(new_n355_), .B2(new_n357_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363_));
  INV_X1    g162(.A(G85gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT0), .B(G57gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n358_), .A2(new_n361_), .A3(new_n360_), .A4(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n332_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n329_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n336_), .B2(new_n373_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n343_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n342_), .A2(new_n376_), .A3(KEYINPUT27), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n320_), .A2(new_n349_), .A3(new_n372_), .A4(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n354_), .A2(new_n357_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT102), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n367_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n355_), .B1(G225gat), .B2(G233gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n379_), .B2(new_n367_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n370_), .B(KEYINPUT33), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n368_), .A2(new_n370_), .B1(new_n387_), .B2(new_n337_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n375_), .A2(KEYINPUT32), .A3(new_n341_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n385_), .A2(new_n386_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n312_), .A2(new_n313_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n315_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n378_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G57gat), .B(G64gat), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n395_), .A2(KEYINPUT11), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(KEYINPUT11), .ZN(new_n397_));
  XOR2_X1   g196(.A(G71gat), .B(G78gat), .Z(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n397_), .A2(new_n398_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G231gat), .A2(G233gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(G231gat), .A3(G233gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G1gat), .B(G8gat), .Z(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(G15gat), .A2(G22gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G15gat), .A2(G22gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(G1gat), .B2(G8gat), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n411_), .A2(new_n413_), .A3(KEYINPUT77), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT77), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G15gat), .B(G22gat), .ZN(new_n416_));
  INV_X1    g215(.A(G1gat), .ZN(new_n417_));
  INV_X1    g216(.A(G8gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT14), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n408_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT77), .B1(new_n411_), .B2(new_n413_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n416_), .A2(new_n415_), .A3(new_n419_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n407_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n406_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n404_), .A2(new_n424_), .A3(new_n405_), .A4(new_n421_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT81), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G127gat), .B(G155gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT80), .ZN(new_n431_));
  XOR2_X1   g230(.A(G183gat), .B(G211gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT17), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n436_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n426_), .A2(new_n427_), .A3(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n429_), .A2(new_n438_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT78), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n428_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n426_), .A2(new_n427_), .A3(KEYINPUT78), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n437_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n394_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G120gat), .B(G148gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(G204gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT5), .B(G176gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT68), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G230gat), .A2(G233gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT66), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT66), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT6), .ZN(new_n462_));
  AND2_X1   g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n460_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n463_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n466_));
  INV_X1    g265(.A(G99gat), .ZN(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n464_), .A2(new_n465_), .A3(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G85gat), .B(G92gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n458_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n464_), .A2(new_n465_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n473_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT9), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT65), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n478_), .A2(new_n364_), .A3(KEYINPUT9), .ZN(new_n479_));
  NOR2_X1   g278(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(G92gat), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT10), .B(G99gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT64), .B(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n475_), .A2(new_n477_), .A3(new_n481_), .A4(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n460_), .A2(new_n462_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n463_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n460_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(KEYINPUT8), .B(new_n476_), .C1(new_n490_), .C2(new_n471_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n474_), .A2(new_n401_), .A3(new_n485_), .A4(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n492_), .A2(KEYINPUT67), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(KEYINPUT67), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n474_), .A2(new_n485_), .A3(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n402_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n457_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n492_), .A2(new_n457_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(KEYINPUT12), .A3(new_n402_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n456_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n493_), .A2(new_n494_), .B1(new_n402_), .B2(new_n496_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n503_), .B(new_n455_), .C1(new_n506_), .C2(new_n457_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(KEYINPUT13), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT13), .B1(new_n505_), .B2(new_n507_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G36gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(G29gat), .ZN(new_n516_));
  INV_X1    g315(.A(G29gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G36gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT69), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT69), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT70), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G29gat), .B(G36gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n514_), .B1(new_n521_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n527_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n519_), .A2(new_n520_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n513_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n422_), .A2(new_n407_), .A3(new_n423_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n407_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n530_), .A2(new_n531_), .A3(new_n513_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n513_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n540_));
  OAI22_X1  g339(.A1(new_n537_), .A2(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n421_), .A2(new_n529_), .A3(new_n424_), .A4(new_n532_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n536_), .B1(new_n543_), .B2(new_n535_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT82), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n546_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT82), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n534_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n550_), .B(new_n545_), .C1(new_n551_), .C2(new_n536_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n547_), .A2(new_n549_), .A3(new_n552_), .A4(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT83), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n547_), .A2(new_n549_), .A3(new_n552_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n555_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n559_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n512_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT72), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n496_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n533_), .B1(new_n496_), .B2(new_n535_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT34), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n496_), .A2(new_n535_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n533_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n496_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT35), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n565_), .B(new_n570_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n572_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT35), .B1(new_n572_), .B2(new_n580_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT75), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(G218gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT73), .B(G190gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT36), .Z(new_n588_));
  AOI21_X1  g387(.A(new_n570_), .B1(new_n577_), .B2(new_n565_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n580_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n578_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n572_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT75), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n583_), .A2(new_n588_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n587_), .A2(KEYINPUT36), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n597_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT76), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT76), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n595_), .A2(new_n601_), .A3(new_n596_), .A4(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n591_), .A2(new_n592_), .A3(new_n588_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(KEYINPUT74), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n596_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n598_), .A2(KEYINPUT74), .A3(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n449_), .A2(new_n564_), .A3(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n610_), .A2(G1gat), .A3(new_n372_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT38), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n595_), .A2(new_n598_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n449_), .A2(new_n564_), .A3(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n372_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(G1324gat));
  NAND2_X1  g415(.A1(new_n349_), .A2(new_n377_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n610_), .A2(G8gat), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT104), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n394_), .A2(new_n448_), .A3(new_n564_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n613_), .ZN(new_n622_));
  OR4_X1    g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n618_), .A4(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n620_), .B1(new_n614_), .B2(new_n618_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n624_), .A3(G8gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n623_), .A2(new_n624_), .A3(new_n627_), .A4(G8gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n619_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n629_), .B(new_n631_), .ZN(G1325gat));
  OAI21_X1  g431(.A(G15gat), .B1(new_n614_), .B2(new_n315_), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n315_), .A2(G15gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n635_), .B1(new_n610_), .B2(new_n636_), .ZN(G1326gat));
  OAI21_X1  g436(.A(G22gat), .B1(new_n614_), .B2(new_n392_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n392_), .A2(G22gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT107), .Z(new_n641_));
  OAI21_X1  g440(.A(new_n639_), .B1(new_n610_), .B2(new_n641_), .ZN(G1327gat));
  NOR3_X1   g441(.A1(new_n512_), .A2(new_n448_), .A3(new_n563_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n394_), .A2(new_n622_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(G29gat), .B1(new_n645_), .B2(new_n371_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n600_), .A2(new_n602_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n394_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT43), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n394_), .A2(new_n650_), .A3(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n643_), .B(KEYINPUT108), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT44), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  AOI211_X1 g455(.A(new_n656_), .B(new_n653_), .C1(new_n649_), .C2(new_n651_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n372_), .A2(new_n517_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n646_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n617_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G36gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n645_), .A2(new_n515_), .A3(new_n617_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT45), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(KEYINPUT46), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  NAND2_X1  g468(.A1(new_n652_), .A2(new_n654_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n656_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n652_), .A2(KEYINPUT44), .A3(new_n654_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n671_), .A2(G43gat), .A3(new_n260_), .A4(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT109), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT109), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n658_), .A2(new_n675_), .A3(G43gat), .A4(new_n260_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n677_), .A2(G43gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(G43gat), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n678_), .B(new_n679_), .C1(new_n644_), .C2(new_n315_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT111), .Z(new_n681_));
  NAND3_X1  g480(.A1(new_n674_), .A2(new_n676_), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT47), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n674_), .A2(new_n676_), .A3(new_n684_), .A4(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1330gat));
  AOI21_X1  g485(.A(G50gat), .B1(new_n645_), .B2(new_n391_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n392_), .A2(new_n299_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n658_), .B2(new_n688_), .ZN(G1331gat));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n511_), .A2(new_n562_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n449_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n692_), .B2(new_n647_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n449_), .A2(KEYINPUT112), .A3(new_n609_), .A4(new_n691_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n692_), .A2(new_n622_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT113), .B1(new_n372_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n696_), .A2(new_n371_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n700_), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n701_), .A2(new_n698_), .B1(KEYINPUT113), .B2(new_n702_), .ZN(G1332gat));
  INV_X1    g502(.A(G64gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n697_), .B2(new_n617_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n705_), .A2(new_n706_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n617_), .A2(new_n704_), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n708_), .A2(new_n709_), .B1(new_n695_), .B2(new_n710_), .ZN(G1333gat));
  INV_X1    g510(.A(G71gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n697_), .B2(new_n260_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT49), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n696_), .A2(new_n712_), .A3(new_n260_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1334gat));
  INV_X1    g515(.A(G78gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n697_), .B2(new_n391_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n718_), .A2(new_n719_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n391_), .A2(new_n717_), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n721_), .A2(new_n722_), .B1(new_n695_), .B2(new_n723_), .ZN(G1335gat));
  NOR3_X1   g523(.A1(new_n511_), .A2(new_n562_), .A3(new_n448_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n394_), .A2(new_n622_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G85gat), .B1(new_n727_), .B2(new_n371_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n652_), .A2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT114), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n652_), .A2(new_n731_), .A3(new_n725_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n478_), .A2(new_n364_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n371_), .B1(new_n480_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT115), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n728_), .B1(new_n733_), .B2(new_n736_), .ZN(G1336gat));
  AOI21_X1  g536(.A(G92gat), .B1(new_n727_), .B2(new_n617_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n617_), .A2(G92gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n733_), .B2(new_n739_), .ZN(G1337gat));
  NAND3_X1  g539(.A1(new_n730_), .A2(new_n260_), .A3(new_n732_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G99gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n727_), .A2(new_n260_), .A3(new_n482_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g544(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n652_), .A2(new_n391_), .A3(new_n725_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G106gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT52), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n727_), .A2(new_n391_), .A3(new_n483_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n748_), .A2(KEYINPUT52), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n747_), .B2(G106gat), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n750_), .B(new_n746_), .C1(new_n752_), .C2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n751_), .A2(new_n756_), .ZN(G1339gat));
  INV_X1    g556(.A(KEYINPUT120), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n618_), .A2(new_n371_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n492_), .A2(KEYINPUT67), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n492_), .A2(KEYINPUT67), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n500_), .B(new_n502_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  INV_X1    g562(.A(new_n457_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n503_), .A2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT55), .A4(new_n502_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n763_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n765_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n453_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n548_), .A2(new_n545_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n555_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n557_), .A2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n503_), .B(new_n453_), .C1(new_n506_), .C2(new_n457_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n762_), .A2(new_n764_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT118), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n767_), .A4(new_n768_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n454_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n772_), .A2(new_n775_), .A3(new_n776_), .A4(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n771_), .A2(KEYINPUT56), .A3(new_n453_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n781_), .B1(new_n780_), .B2(new_n454_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n775_), .A4(new_n776_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n603_), .A2(new_n608_), .A3(new_n785_), .A4(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n772_), .A2(new_n562_), .A3(new_n776_), .A4(new_n782_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n505_), .A2(new_n507_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n775_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n613_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n613_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n790_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n447_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n509_), .A2(new_n510_), .A3(new_n447_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n563_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT13), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n792_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n448_), .A3(new_n508_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n806_), .A2(new_n562_), .A3(KEYINPUT117), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n803_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n609_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n803_), .A2(new_n807_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT54), .B1(new_n647_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n759_), .B1(new_n800_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n314_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT59), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n799_), .A2(new_n447_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  NOR4_X1   g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n314_), .A4(new_n759_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n758_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n759_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n810_), .A2(new_n812_), .ZN(new_n822_));
  AOI221_X4 g621(.A(new_n796_), .B1(new_n598_), .B2(new_n595_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT57), .B1(new_n794_), .B2(new_n613_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n448_), .B1(new_n825_), .B2(new_n790_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n815_), .B(new_n821_), .C1(new_n822_), .C2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n818_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n814_), .A2(KEYINPUT59), .A3(new_n815_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(KEYINPUT120), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n820_), .A2(G113gat), .A3(new_n830_), .A4(new_n562_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n827_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n562_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n833_), .A2(KEYINPUT119), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(KEYINPUT119), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n831_), .A2(new_n834_), .A3(new_n835_), .ZN(G1340gat));
  NOR2_X1   g635(.A1(new_n511_), .A2(G120gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n832_), .B1(KEYINPUT60), .B2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n512_), .C1(new_n816_), .C2(new_n819_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(KEYINPUT60), .B2(new_n838_), .ZN(G1341gat));
  INV_X1    g640(.A(G127gat), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n447_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n820_), .A2(new_n830_), .A3(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n827_), .B2(new_n447_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n844_), .A2(KEYINPUT121), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT121), .B1(new_n844_), .B2(new_n845_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1342gat));
  AND4_X1   g647(.A1(G134gat), .A2(new_n820_), .A3(new_n647_), .A4(new_n830_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G134gat), .B1(new_n832_), .B2(new_n622_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1343gat));
  NOR3_X1   g650(.A1(new_n817_), .A2(new_n319_), .A3(new_n759_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n562_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n512_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g655(.A1(new_n852_), .A2(new_n448_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n857_), .B(new_n860_), .ZN(G1346gat));
  AOI21_X1  g660(.A(G162gat), .B1(new_n852_), .B2(new_n622_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n647_), .A2(G162gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n852_), .B2(new_n863_), .ZN(G1347gat));
  AOI21_X1  g663(.A(new_n371_), .B1(new_n800_), .B2(new_n813_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(new_n617_), .A3(new_n815_), .A4(new_n562_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G169gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n868_));
  INV_X1    g667(.A(new_n219_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n867_), .B(new_n868_), .C1(new_n869_), .C2(new_n866_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  INV_X1    g670(.A(new_n868_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n866_), .A2(G169gat), .A3(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n871_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n871_), .B1(new_n870_), .B2(new_n873_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1348gat));
  OAI211_X1 g676(.A(new_n372_), .B(new_n617_), .C1(new_n822_), .C2(new_n826_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n314_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n512_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n448_), .ZN(new_n882_));
  MUX2_X1   g681(.A(new_n324_), .B(G183gat), .S(new_n882_), .Z(G1350gat));
  INV_X1    g682(.A(new_n879_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G190gat), .B1(new_n884_), .B2(new_n609_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n879_), .A2(new_n233_), .A3(new_n622_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1351gat));
  OAI21_X1  g686(.A(KEYINPUT126), .B1(new_n878_), .B2(new_n319_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889_));
  INV_X1    g688(.A(new_n319_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n865_), .A2(new_n889_), .A3(new_n617_), .A4(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n562_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n512_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n892_), .B2(new_n448_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT63), .B(G211gat), .Z(new_n899_));
  AOI211_X1 g698(.A(new_n447_), .B(new_n899_), .C1(new_n888_), .C2(new_n891_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT127), .B1(new_n898_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n899_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n892_), .A2(new_n448_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n447_), .B1(new_n888_), .B2(new_n891_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n903_), .B(new_n904_), .C1(new_n905_), .C2(new_n897_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n901_), .A2(new_n906_), .ZN(G1354gat));
  AOI21_X1  g706(.A(G218gat), .B1(new_n892_), .B2(new_n622_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n609_), .B1(new_n888_), .B2(new_n891_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(G218gat), .B2(new_n909_), .ZN(G1355gat));
endmodule


