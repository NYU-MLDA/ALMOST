//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n941_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n987_, new_n988_, new_n990_, new_n991_,
    new_n992_, new_n994_, new_n995_, new_n996_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1003_, new_n1004_, new_n1005_, new_n1006_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT8), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT66), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n202_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n205_), .B1(new_n210_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n203_), .A2(KEYINPUT66), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n213_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT9), .A3(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(KEYINPUT65), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G92gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n223_), .A2(KEYINPUT9), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n232_), .A2(new_n233_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n217_), .A2(new_n219_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n225_), .B(new_n226_), .C1(KEYINPUT66), .C2(new_n203_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n216_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n207_), .A2(new_n209_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n218_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G43gat), .B(G50gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n245_), .A2(KEYINPUT15), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT15), .B1(new_n245_), .B2(new_n247_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G232gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT34), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(KEYINPUT35), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n245_), .A2(new_n247_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n235_), .A2(new_n255_), .A3(new_n240_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT35), .A3(new_n253_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(KEYINPUT35), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n251_), .A2(new_n259_), .A3(new_n254_), .A4(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G190gat), .B(G218gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G134gat), .B(G162gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT36), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n258_), .A2(new_n265_), .A3(new_n260_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(KEYINPUT36), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT37), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n269_), .A2(KEYINPUT37), .A3(new_n270_), .A4(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G127gat), .B(G155gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G183gat), .B(G211gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n282_), .A2(KEYINPUT17), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(KEYINPUT17), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT73), .ZN(new_n285_));
  XOR2_X1   g084(.A(G1gat), .B(G8gat), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(G15gat), .A2(G22gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G15gat), .A2(G22gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT14), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(G1gat), .B2(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT70), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G22gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n296_));
  INV_X1    g095(.A(G1gat), .ZN(new_n297_));
  INV_X1    g096(.A(G8gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT14), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n293_), .A2(new_n294_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n294_), .B1(new_n293_), .B2(new_n300_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n287_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n290_), .A2(new_n292_), .A3(KEYINPUT70), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n296_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT71), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n293_), .A2(new_n294_), .A3(new_n300_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n286_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G64gat), .ZN(new_n314_));
  INV_X1    g113(.A(G78gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G71gat), .ZN(new_n316_));
  INV_X1    g115(.A(G71gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G78gat), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n314_), .A2(KEYINPUT11), .A3(new_n316_), .A4(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G64gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G57gat), .ZN(new_n321_));
  INV_X1    g120(.A(G57gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G64gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n323_), .A3(KEYINPUT11), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n318_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n314_), .A2(KEYINPUT11), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n313_), .B(new_n319_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(new_n323_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n313_), .B1(new_n333_), .B2(new_n319_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n311_), .B(new_n312_), .C1(new_n329_), .C2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n319_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT67), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n309_), .A2(new_n310_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n309_), .A2(new_n310_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n328_), .B(new_n337_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT73), .B1(new_n283_), .B2(new_n284_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n285_), .A2(new_n335_), .A3(new_n340_), .A4(new_n341_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n319_), .B(new_n333_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n311_), .A2(new_n336_), .A3(new_n312_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n283_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT74), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n232_), .A2(new_n233_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n348_), .A2(new_n238_), .A3(new_n227_), .A4(new_n222_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(new_n239_), .B2(new_n218_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n217_), .A2(new_n219_), .ZN(new_n351_));
  OAI22_X1  g150(.A1(new_n350_), .A2(new_n351_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT12), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n333_), .A2(KEYINPUT12), .A3(new_n319_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n352_), .A2(new_n353_), .B1(new_n241_), .B2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n235_), .A2(new_n337_), .A3(new_n328_), .A4(new_n240_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G230gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT64), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n357_), .A2(KEYINPUT68), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT68), .B1(new_n357_), .B2(new_n359_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n356_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n352_), .A2(new_n357_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G120gat), .B(G148gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT5), .ZN(new_n368_));
  XOR2_X1   g167(.A(G176gat), .B(G204gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n366_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT13), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n372_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n277_), .A2(new_n347_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT26), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G190gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT79), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(G183gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(new_n377_), .A3(G190gat), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n379_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT78), .B(G190gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT26), .ZN(new_n387_));
  INV_X1    g186(.A(G183gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(KEYINPUT25), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n381_), .A2(G183gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(KEYINPUT77), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n385_), .A2(new_n387_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT24), .ZN(new_n393_));
  INV_X1    g192(.A(G169gat), .ZN(new_n394_));
  INV_X1    g193(.A(G176gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT23), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT80), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n396_), .A2(new_n399_), .A3(new_n403_), .A4(new_n400_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n394_), .A2(new_n395_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n392_), .A2(new_n405_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT81), .B1(new_n394_), .B2(KEYINPUT22), .ZN(new_n411_));
  AOI21_X1  g210(.A(G176gat), .B1(new_n394_), .B2(KEYINPUT22), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT22), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(G169gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n406_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT82), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n420_), .A3(new_n417_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n386_), .A2(new_n388_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n399_), .A2(new_n400_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n419_), .A2(new_n421_), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n410_), .A2(new_n425_), .A3(KEYINPUT30), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT30), .B1(new_n410_), .B2(new_n425_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n376_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n410_), .A2(new_n425_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n376_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(G15gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G43gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n429_), .A2(new_n434_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n439_), .B1(new_n429_), .B2(new_n434_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G127gat), .B(G134gat), .Z(new_n443_));
  XOR2_X1   g242(.A(G113gat), .B(G120gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT31), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT84), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n441_), .A2(new_n442_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n446_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n429_), .A2(new_n434_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n438_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n453_), .B1(new_n455_), .B2(new_n440_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n451_), .A2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(G141gat), .A2(G148gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT2), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G141gat), .A2(G148gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT3), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G141gat), .A2(G148gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT2), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n459_), .A2(new_n462_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(G155gat), .A2(G162gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(G155gat), .A2(G162gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT1), .ZN(new_n472_));
  INV_X1    g271(.A(G141gat), .ZN(new_n473_));
  INV_X1    g272(.A(G148gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n463_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n472_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AND3_X1   g278(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n480_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n481_));
  OR2_X1    g280(.A1(G155gat), .A2(G162gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT1), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G155gat), .A2(G162gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT85), .B1(new_n481_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n471_), .B1(new_n479_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT28), .B1(new_n487_), .B2(KEYINPUT29), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n478_), .B1(new_n472_), .B2(new_n477_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n458_), .A2(new_n460_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n485_), .A2(new_n490_), .A3(KEYINPUT85), .A4(new_n476_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n489_), .A2(new_n491_), .B1(new_n470_), .B2(new_n467_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT28), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT29), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n487_), .A2(KEYINPUT29), .ZN(new_n497_));
  INV_X1    g296(.A(G218gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G211gat), .ZN(new_n499_));
  INV_X1    g298(.A(G211gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G218gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT89), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G211gat), .B(G218gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G197gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G204gat), .ZN(new_n508_));
  INV_X1    g307(.A(G204gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(G197gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n503_), .A2(new_n506_), .A3(KEYINPUT21), .A4(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G197gat), .B(G204gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n502_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(KEYINPUT21), .A3(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n515_), .A2(KEYINPUT88), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT88), .B1(new_n515_), .B2(new_n519_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n512_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n496_), .A2(new_n497_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n497_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(new_n488_), .A3(new_n495_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G228gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(new_n315_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n213_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G22gat), .B(G50gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n523_), .A2(new_n525_), .A3(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G1gat), .B(G29gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G57gat), .B(G85gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n443_), .B(new_n444_), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n487_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n492_), .A2(new_n445_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(KEYINPUT4), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G225gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  OR3_X1    g345(.A1(new_n492_), .A2(KEYINPUT4), .A3(new_n445_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n544_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n542_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n540_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n549_), .A3(new_n540_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  AOI211_X1 g353(.A(new_n552_), .B(new_n540_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n535_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n457_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT27), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G226gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT19), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT90), .Z(new_n562_));
  AND4_X1   g361(.A1(KEYINPUT21), .A2(new_n503_), .A3(new_n506_), .A4(new_n511_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n518_), .A2(KEYINPUT21), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n516_), .B2(new_n513_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT21), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT87), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT87), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT21), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n504_), .B1(new_n511_), .B2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n564_), .B1(new_n566_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n515_), .A2(new_n519_), .A3(KEYINPUT88), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n563_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(G190gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n388_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n399_), .A2(new_n400_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT22), .B(G169gat), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n406_), .B1(new_n581_), .B2(new_n395_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n401_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n390_), .A2(new_n389_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT26), .B(G190gat), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n408_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n580_), .A2(new_n582_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT92), .B1(new_n575_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n578_), .A2(new_n579_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n578_), .A2(new_n579_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n582_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n586_), .A2(new_n583_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n522_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT20), .B1(new_n430_), .B2(new_n522_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n562_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT20), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n575_), .B2(new_n587_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n561_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n410_), .A2(new_n425_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n600_), .B(new_n601_), .C1(new_n575_), .C2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G8gat), .B(G36gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G64gat), .B(G92gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n598_), .A2(new_n603_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n598_), .B2(new_n603_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n559_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n598_), .A2(new_n603_), .A3(new_n608_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n599_), .B1(new_n602_), .B2(new_n575_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n562_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(new_n588_), .A4(new_n595_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n602_), .A2(new_n575_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT20), .B1(new_n522_), .B2(new_n594_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n561_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n612_), .B(KEYINPUT27), .C1(new_n619_), .C2(new_n608_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n611_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n558_), .A2(new_n621_), .A3(KEYINPUT98), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n457_), .A2(new_n557_), .A3(new_n611_), .A4(new_n620_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n554_), .A2(new_n556_), .ZN(new_n627_));
  AND4_X1   g426(.A1(new_n627_), .A2(new_n611_), .A3(new_n535_), .A4(new_n620_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n609_), .A2(new_n610_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n553_), .A2(KEYINPUT33), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n548_), .A2(new_n631_), .A3(new_n549_), .A4(new_n540_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n544_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n540_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT95), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n544_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n639_), .A2(new_n640_), .A3(new_n636_), .A4(new_n635_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n629_), .A2(KEYINPUT96), .A3(new_n633_), .A4(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n598_), .A2(new_n603_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n608_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n646_), .A2(new_n633_), .A3(new_n612_), .A4(new_n642_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n553_), .A2(new_n552_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n550_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n555_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n608_), .A2(KEYINPUT32), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n598_), .A2(new_n603_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(new_n653_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n643_), .A2(new_n649_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n535_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n628_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n626_), .B1(new_n660_), .B2(new_n457_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(G113gat), .B(G141gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(G169gat), .B(G197gat), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n662_), .B(new_n663_), .Z(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n303_), .A2(new_n250_), .A3(new_n308_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(G229gat), .A2(G233gat), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT76), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT75), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n309_), .B2(new_n255_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n255_), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT75), .B(new_n672_), .C1(new_n303_), .C2(new_n308_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n668_), .B(new_n669_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n309_), .A2(new_n255_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n308_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n286_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n255_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT75), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n309_), .A2(new_n670_), .A3(new_n255_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n674_), .B1(new_n681_), .B2(new_n667_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n680_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n669_), .B1(new_n683_), .B2(new_n668_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n665_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n667_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n671_), .A2(new_n673_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(new_n675_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n668_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT76), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n688_), .A2(new_n690_), .A3(new_n674_), .A4(new_n664_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n685_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n661_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n661_), .A2(KEYINPUT99), .A3(new_n692_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n375_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n627_), .A2(G1gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT38), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(KEYINPUT38), .A3(new_n698_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n271_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n347_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n457_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n648_), .A2(new_n647_), .B1(new_n652_), .B2(new_n656_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n535_), .B1(new_n706_), .B2(new_n643_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n707_), .B2(new_n628_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n704_), .B1(new_n708_), .B2(new_n626_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n373_), .A2(new_n374_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(new_n692_), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G1gat), .B1(new_n712_), .B2(new_n627_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n701_), .A2(new_n702_), .A3(new_n713_), .ZN(G1324gat));
  INV_X1    g513(.A(new_n621_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n697_), .A2(new_n298_), .A3(new_n715_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n712_), .A2(KEYINPUT100), .A3(new_n621_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n298_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT39), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT100), .B1(new_n712_), .B2(new_n621_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n716_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n716_), .B(new_n724_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1325gat));
  OAI21_X1  g527(.A(G15gat), .B1(new_n712_), .B2(new_n705_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n730_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n697_), .A2(new_n436_), .A3(new_n457_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(G1326gat));
  OAI21_X1  g533(.A(G22gat), .B1(new_n712_), .B2(new_n659_), .ZN(new_n735_));
  XOR2_X1   g534(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n659_), .A2(G22gat), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT104), .Z(new_n739_));
  NAND2_X1  g538(.A1(new_n697_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(G1327gat));
  NAND2_X1  g540(.A1(new_n695_), .A2(new_n696_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n347_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n271_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(new_n710_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n627_), .A2(G29gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n692_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n710_), .A2(new_n748_), .A3(new_n347_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT43), .B(new_n277_), .C1(new_n708_), .C2(new_n626_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n751_));
  INV_X1    g550(.A(new_n277_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n661_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT44), .B(new_n749_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n652_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(G29gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G29gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n747_), .B1(new_n761_), .B2(new_n762_), .ZN(G1328gat));
  NAND3_X1  g562(.A1(new_n756_), .A2(new_n715_), .A3(new_n757_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G36gat), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n621_), .A2(G36gat), .ZN(new_n766_));
  INV_X1    g565(.A(new_n696_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT99), .B1(new_n661_), .B2(new_n692_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n745_), .B(new_n766_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT106), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n742_), .A2(new_n772_), .A3(new_n745_), .A4(new_n766_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n770_), .A2(new_n771_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n765_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT46), .B(new_n765_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1329gat));
  XNOR2_X1  g579(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(G43gat), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n705_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n756_), .A2(new_n757_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n742_), .A2(new_n457_), .A3(new_n745_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n783_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n785_), .A2(new_n786_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n786_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n782_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n785_), .A2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT108), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n785_), .A2(new_n786_), .A3(new_n788_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n781_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1330gat));
  INV_X1    g595(.A(G50gat), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n659_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n742_), .A2(new_n535_), .A3(new_n745_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n758_), .A2(new_n798_), .B1(new_n797_), .B2(new_n799_), .ZN(G1331gat));
  NOR2_X1   g599(.A1(new_n711_), .A2(new_n692_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n709_), .A2(new_n801_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n802_), .A2(new_n322_), .A3(new_n627_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT110), .Z(new_n804_));
  AOI21_X1  g603(.A(new_n692_), .B1(new_n708_), .B2(new_n626_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n277_), .A2(new_n347_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n710_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n808_), .A2(KEYINPUT109), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(KEYINPUT109), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n652_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n804_), .B1(new_n322_), .B2(new_n811_), .ZN(G1332gat));
  OAI21_X1  g611(.A(G64gat), .B1(new_n802_), .B2(new_n621_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT48), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n808_), .A2(new_n320_), .A3(new_n715_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1333gat));
  OAI21_X1  g615(.A(G71gat), .B1(new_n802_), .B2(new_n705_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT49), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n808_), .A2(new_n317_), .A3(new_n457_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1334gat));
  OAI21_X1  g619(.A(G78gat), .B1(new_n802_), .B2(new_n659_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT50), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n808_), .A2(new_n315_), .A3(new_n535_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1335gat));
  OR2_X1    g623(.A1(new_n750_), .A2(new_n753_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n711_), .A2(new_n692_), .A3(new_n347_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G85gat), .B1(new_n827_), .B2(new_n627_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n744_), .A2(new_n711_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n805_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n223_), .A3(new_n652_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(G1336gat));
  AOI21_X1  g632(.A(G92gat), .B1(new_n831_), .B2(new_n715_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n827_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n621_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(G1337gat));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT51), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n457_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n830_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n835_), .A2(new_n457_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(G99gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n838_), .A2(KEYINPUT51), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1338gat));
  NAND3_X1  g644(.A1(new_n831_), .A2(new_n213_), .A3(new_n535_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n825_), .A2(new_n535_), .A3(new_n826_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(KEYINPUT52), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n213_), .B1(new_n848_), .B2(KEYINPUT52), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n847_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n846_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT53), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n855_), .B(new_n846_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1339gat));
  NOR2_X1   g656(.A1(new_n715_), .A2(new_n627_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n705_), .A2(new_n535_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n366_), .A2(new_n370_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n241_), .A2(new_n355_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n240_), .A2(new_n235_), .B1(new_n337_), .B2(new_n328_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n862_), .B(new_n357_), .C1(new_n863_), .C2(KEYINPUT12), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n352_), .A2(new_n353_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n867_), .A2(KEYINPUT113), .A3(new_n357_), .A4(new_n862_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n868_), .A3(new_n364_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n362_), .A2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n356_), .B(KEYINPUT55), .C1(new_n360_), .C2(new_n361_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n873_), .A2(KEYINPUT56), .A3(new_n370_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n873_), .B2(new_n370_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n692_), .B(new_n861_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n683_), .A2(new_n686_), .A3(new_n666_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n877_), .B(new_n665_), .C1(new_n686_), .C2(new_n681_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n371_), .A2(new_n691_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(KEYINPUT57), .A3(new_n703_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n691_), .A2(new_n861_), .A3(new_n878_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT58), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n884_), .B(new_n887_), .C1(new_n875_), .C2(new_n874_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n752_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n880_), .A2(new_n703_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n271_), .B1(new_n876_), .B2(new_n879_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n883_), .A2(new_n890_), .A3(new_n893_), .A4(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n743_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n806_), .A2(new_n711_), .A3(new_n898_), .A4(new_n748_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT54), .B1(new_n375_), .B2(new_n692_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n860_), .B1(new_n897_), .B2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(KEYINPUT59), .ZN(new_n903_));
  INV_X1    g702(.A(new_n901_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n896_), .B2(new_n743_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n905_), .A2(new_n906_), .A3(new_n860_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n903_), .A2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G113gat), .B1(new_n908_), .B2(new_n748_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n902_), .ZN(new_n910_));
  OR3_X1    g709(.A1(new_n910_), .A2(G113gat), .A3(new_n748_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1340gat));
  OAI21_X1  g711(.A(G120gat), .B1(new_n908_), .B2(new_n711_), .ZN(new_n913_));
  INV_X1    g712(.A(G120gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT116), .B1(new_n914_), .B2(KEYINPUT60), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n711_), .B2(KEYINPUT60), .ZN(new_n916_));
  MUX2_X1   g715(.A(KEYINPUT116), .B(new_n915_), .S(new_n916_), .Z(new_n917_));
  OAI21_X1  g716(.A(new_n913_), .B1(new_n910_), .B2(new_n917_), .ZN(G1341gat));
  INV_X1    g717(.A(G127gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n743_), .A2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n903_), .B2(new_n907_), .ZN(new_n921_));
  AOI211_X1 g720(.A(KEYINPUT117), .B(G127gat), .C1(new_n902_), .C2(new_n347_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n897_), .A2(new_n901_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n860_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n924_), .A2(new_n347_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n923_), .B1(new_n926_), .B2(new_n919_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n921_), .B1(new_n922_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n921_), .B(KEYINPUT118), .C1(new_n927_), .C2(new_n922_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1342gat));
  AOI21_X1  g731(.A(G134gat), .B1(new_n902_), .B2(new_n271_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n908_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n752_), .A2(G134gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT119), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n933_), .B1(new_n934_), .B2(new_n936_), .ZN(G1343gat));
  NAND4_X1  g736(.A1(new_n924_), .A2(new_n535_), .A3(new_n705_), .A4(new_n858_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n748_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(new_n473_), .ZN(G1344gat));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n711_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n474_), .ZN(G1345gat));
  NOR2_X1   g741(.A1(new_n938_), .A2(new_n743_), .ZN(new_n943_));
  XOR2_X1   g742(.A(KEYINPUT61), .B(G155gat), .Z(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n938_), .B2(new_n277_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n703_), .A2(G162gat), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n938_), .B2(new_n947_), .ZN(G1347gat));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949_));
  AOI21_X1  g748(.A(KEYINPUT115), .B1(new_n894_), .B2(KEYINPUT57), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n277_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n892_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n952_), .B1(new_n880_), .B2(new_n703_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n950_), .A2(new_n951_), .A3(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n347_), .B1(new_n954_), .B2(new_n895_), .ZN(new_n955_));
  OAI211_X1 g754(.A(new_n715_), .B(new_n558_), .C1(new_n955_), .C2(new_n904_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n692_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n949_), .B1(new_n958_), .B2(G169gat), .ZN(new_n959_));
  AOI211_X1 g758(.A(KEYINPUT62), .B(new_n394_), .C1(new_n957_), .C2(new_n692_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n621_), .B1(new_n897_), .B2(new_n901_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n961_), .B1(new_n962_), .B2(new_n558_), .ZN(new_n963_));
  INV_X1    g762(.A(new_n558_), .ZN(new_n964_));
  NOR4_X1   g763(.A1(new_n905_), .A2(KEYINPUT120), .A3(new_n621_), .A4(new_n964_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n963_), .A2(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n692_), .A2(new_n581_), .ZN(new_n967_));
  OAI22_X1  g766(.A1(new_n959_), .A2(new_n960_), .B1(new_n966_), .B2(new_n967_), .ZN(G1348gat));
  NOR3_X1   g767(.A1(new_n956_), .A2(new_n395_), .A3(new_n711_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n956_), .A2(KEYINPUT120), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n962_), .A2(new_n961_), .A3(new_n558_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n711_), .B1(new_n970_), .B2(new_n971_), .ZN(new_n972_));
  OAI21_X1  g771(.A(KEYINPUT121), .B1(new_n972_), .B2(G176gat), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT121), .ZN(new_n974_));
  OAI211_X1 g773(.A(new_n974_), .B(new_n395_), .C1(new_n966_), .C2(new_n711_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n969_), .B1(new_n973_), .B2(new_n975_), .ZN(G1349gat));
  NOR2_X1   g775(.A1(new_n743_), .A2(new_n584_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n977_), .B1(new_n963_), .B2(new_n965_), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n978_), .A2(new_n979_), .ZN(new_n980_));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n957_), .A2(new_n981_), .A3(new_n347_), .ZN(new_n982_));
  OAI21_X1  g781(.A(KEYINPUT123), .B1(new_n956_), .B2(new_n743_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n982_), .A2(new_n388_), .A3(new_n983_), .ZN(new_n984_));
  OAI211_X1 g783(.A(KEYINPUT122), .B(new_n977_), .C1(new_n963_), .C2(new_n965_), .ZN(new_n985_));
  AND3_X1   g784(.A1(new_n980_), .A2(new_n984_), .A3(new_n985_), .ZN(G1350gat));
  OAI21_X1  g785(.A(G190gat), .B1(new_n966_), .B2(new_n277_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n271_), .A2(new_n585_), .ZN(new_n988_));
  OAI21_X1  g787(.A(new_n987_), .B1(new_n966_), .B2(new_n988_), .ZN(G1351gat));
  NOR3_X1   g788(.A1(new_n457_), .A2(new_n652_), .A3(new_n659_), .ZN(new_n990_));
  AND2_X1   g789(.A1(new_n962_), .A2(new_n990_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n991_), .A2(new_n692_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n992_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g792(.A1(new_n991_), .A2(new_n710_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n995_));
  XOR2_X1   g794(.A(new_n995_), .B(KEYINPUT125), .Z(new_n996_));
  XNOR2_X1  g795(.A(new_n994_), .B(new_n996_), .ZN(G1353gat));
  NAND2_X1  g796(.A1(new_n991_), .A2(new_n347_), .ZN(new_n998_));
  NOR2_X1   g797(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n999_));
  AND2_X1   g798(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1000_));
  NOR3_X1   g799(.A1(new_n998_), .A2(new_n999_), .A3(new_n1000_), .ZN(new_n1001_));
  AOI21_X1  g800(.A(new_n1001_), .B1(new_n998_), .B2(new_n999_), .ZN(G1354gat));
  NAND3_X1  g801(.A1(new_n962_), .A2(new_n271_), .A3(new_n990_), .ZN(new_n1003_));
  XNOR2_X1  g802(.A(new_n1003_), .B(KEYINPUT126), .ZN(new_n1004_));
  XNOR2_X1  g803(.A(KEYINPUT127), .B(G218gat), .ZN(new_n1005_));
  NOR2_X1   g804(.A1(new_n277_), .A2(new_n1005_), .ZN(new_n1006_));
  AOI22_X1  g805(.A1(new_n1004_), .A2(new_n1005_), .B1(new_n991_), .B2(new_n1006_), .ZN(G1355gat));
endmodule


