//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n924_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G218gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G211gat), .ZN(new_n209_));
  INV_X1    g008(.A(G211gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G218gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT21), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G197gat), .B(G204gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT87), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(KEYINPUT87), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n213_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G197gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G204gat), .ZN(new_n219_));
  INV_X1    g018(.A(G204gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G197gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT85), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT21), .B1(new_n219_), .B2(KEYINPUT85), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n221_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n209_), .B(new_n211_), .C1(new_n225_), .C2(KEYINPUT21), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT86), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT21), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n212_), .B1(new_n228_), .B2(new_n214_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT85), .ZN(new_n230_));
  OR3_X1    g029(.A1(new_n220_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT21), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n217_), .B1(new_n227_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(G183gat), .ZN(new_n237_));
  INV_X1    g036(.A(G183gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(KEYINPUT25), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT92), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT26), .B(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(KEYINPUT25), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(G183gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT92), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT24), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(G169gat), .B2(G176gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT77), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(G169gat), .B2(G176gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n246_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT93), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT93), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n246_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n250_), .A2(new_n252_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n247_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n255_), .A2(new_n257_), .A3(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n258_), .B(KEYINPUT23), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(G183gat), .B2(G190gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT78), .B(G176gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT22), .B(G169gat), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n266_), .A2(new_n267_), .B1(G169gat), .B2(G176gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n235_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n214_), .B(KEYINPUT87), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(KEYINPUT21), .A3(new_n212_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n229_), .A2(new_n233_), .A3(new_n232_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n233_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n276_), .A2(new_n253_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n262_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n269_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT20), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT19), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT91), .ZN(new_n283_));
  OR3_X1    g082(.A1(new_n270_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n282_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT20), .ZN(new_n286_));
  INV_X1    g085(.A(new_n269_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n261_), .A2(new_n247_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n264_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n254_), .B2(KEYINPUT93), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n287_), .B1(new_n290_), .B2(new_n257_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n291_), .B2(new_n235_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n277_), .A2(new_n262_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT95), .B1(new_n235_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT95), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n275_), .A2(new_n295_), .A3(new_n279_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n285_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT99), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n284_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AOI211_X1 g099(.A(KEYINPUT99), .B(new_n285_), .C1(new_n292_), .C2(new_n297_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n202_), .B(new_n207_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n283_), .B1(new_n270_), .B2(new_n280_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT94), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OAI211_X1 g104(.A(KEYINPUT94), .B(new_n283_), .C1(new_n270_), .C2(new_n280_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n292_), .A2(new_n297_), .A3(new_n285_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n305_), .A2(new_n206_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n308_), .A2(KEYINPUT27), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n294_), .A2(new_n296_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n263_), .A2(new_n269_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT20), .B1(new_n312_), .B2(new_n275_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n282_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT99), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n298_), .A2(new_n299_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n284_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n202_), .B1(new_n317_), .B2(new_n207_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n207_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n308_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  OAI22_X1  g121(.A1(new_n310_), .A2(new_n318_), .B1(new_n322_), .B2(KEYINPUT27), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G78gat), .B(G106gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n325_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(new_n328_), .B2(new_n327_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n325_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT83), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n326_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT83), .B1(new_n327_), .B2(new_n325_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340_));
  NOR4_X1   g139(.A1(new_n340_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT80), .B1(new_n331_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n333_), .A2(KEYINPUT81), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT81), .B1(new_n333_), .B2(new_n344_), .ZN(new_n346_));
  OAI22_X1  g145(.A1(new_n341_), .A2(new_n343_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT82), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n350_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(KEYINPUT84), .B(new_n339_), .C1(new_n347_), .C2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n353_), .ZN(new_n356_));
  INV_X1    g155(.A(G141gat), .ZN(new_n357_));
  INV_X1    g156(.A(G148gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n342_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n340_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n331_), .A2(KEYINPUT80), .A3(new_n342_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n333_), .A2(new_n344_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n333_), .A2(KEYINPUT81), .A3(new_n344_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n356_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT84), .B1(new_n368_), .B2(new_n339_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n334_), .B1(new_n355_), .B2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n235_), .B1(new_n370_), .B2(KEYINPUT29), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n275_), .B2(KEYINPUT88), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n334_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n339_), .B1(new_n347_), .B2(new_n353_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n376_), .B1(new_n379_), .B2(new_n354_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n275_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(new_n373_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n324_), .B1(new_n375_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n371_), .A2(new_n374_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n373_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n324_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(KEYINPUT89), .A3(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT28), .B1(new_n370_), .B2(KEYINPUT29), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT28), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n380_), .A2(new_n391_), .A3(new_n381_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G22gat), .B(G50gat), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n398_), .B(new_n324_), .C1(new_n375_), .C2(new_n383_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n389_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n384_), .A2(KEYINPUT90), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT90), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n402_), .B(new_n324_), .C1(new_n375_), .C2(new_n383_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n401_), .A2(new_n403_), .A3(new_n396_), .A4(new_n388_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n323_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G127gat), .B(G134gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G113gat), .B(G120gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n334_), .B(new_n412_), .C1(new_n355_), .C2(new_n369_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n412_), .B(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n413_), .B(KEYINPUT4), .C1(new_n380_), .C2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT97), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n379_), .A2(new_n354_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n415_), .B1(new_n418_), .B2(new_n334_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n417_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  NOR4_X1   g221(.A1(new_n380_), .A2(new_n415_), .A3(KEYINPUT97), .A4(new_n420_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n409_), .B(new_n416_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n413_), .B(new_n408_), .C1(new_n380_), .C2(new_n415_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G85gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT0), .B(G57gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n424_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT101), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n416_), .A2(new_n409_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n412_), .B(KEYINPUT79), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n370_), .A2(new_n436_), .A3(new_n421_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT97), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n419_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n431_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT101), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n424_), .A2(new_n425_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n434_), .A2(new_n443_), .B1(new_n444_), .B2(new_n429_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G15gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT30), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n293_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(new_n415_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451_));
  INV_X1    g250(.A(G43gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT31), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n450_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n445_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n407_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT102), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n319_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n434_), .A2(new_n443_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n444_), .A2(new_n429_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT100), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n317_), .B2(new_n460_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n465_), .B(new_n460_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n433_), .A2(KEYINPUT98), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT98), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n441_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n440_), .A2(new_n408_), .A3(new_n416_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n419_), .B1(new_n380_), .B2(new_n412_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n430_), .B1(new_n476_), .B2(new_n409_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n424_), .A2(KEYINPUT33), .A3(new_n432_), .ZN(new_n479_));
  AND4_X1   g278(.A1(new_n308_), .A2(new_n478_), .A3(new_n320_), .A4(new_n479_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n464_), .A2(new_n469_), .B1(new_n474_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n459_), .B1(new_n481_), .B2(new_n405_), .ZN(new_n482_));
  AOI211_X1 g281(.A(KEYINPUT101), .B(new_n431_), .C1(new_n435_), .C2(new_n440_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n442_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n463_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n461_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n460_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT100), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n485_), .A2(new_n486_), .A3(new_n488_), .A4(new_n467_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n478_), .A2(new_n479_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n474_), .A2(new_n322_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n405_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(KEYINPUT102), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n405_), .A2(new_n445_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT104), .B1(new_n323_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n318_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n302_), .A2(new_n309_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT27), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n497_), .A2(new_n498_), .B1(new_n499_), .B2(new_n321_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT104), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n485_), .B1(new_n404_), .B2(new_n400_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n482_), .A2(new_n494_), .A3(new_n496_), .A4(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n458_), .B1(new_n504_), .B2(new_n455_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G29gat), .B(G36gat), .Z(new_n506_));
  XOR2_X1   g305(.A(G43gat), .B(G50gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT15), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  INV_X1    g309(.A(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G8gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n508_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(new_n516_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n518_), .B(new_n516_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G113gat), .B(G141gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT76), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n525_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n505_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT37), .ZN(new_n534_));
  INV_X1    g333(.A(G99gat), .ZN(new_n535_));
  INV_X1    g334(.A(G106gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT6), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT6), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(G99gat), .A3(G106gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT65), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n542_), .A2(KEYINPUT9), .ZN(new_n543_));
  INV_X1    g342(.A(G85gat), .ZN(new_n544_));
  INV_X1    g343(.A(G92gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n542_), .B2(KEYINPUT9), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT10), .B(G99gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT64), .Z(new_n549_));
  OAI221_X1 g348(.A(new_n540_), .B1(new_n543_), .B2(new_n547_), .C1(new_n549_), .C2(G106gat), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT8), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n540_), .B(KEYINPUT66), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT67), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT66), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n540_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT67), .ZN(new_n557_));
  NOR2_X1   g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT7), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n554_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n546_), .A2(new_n541_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n551_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  AOI211_X1 g362(.A(KEYINPUT8), .B(new_n561_), .C1(new_n559_), .C2(new_n540_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n508_), .B(new_n550_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT70), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n550_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n509_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n572_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n569_), .A2(new_n570_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(KEYINPUT70), .A3(new_n509_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n573_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n565_), .A2(new_n571_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n577_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n589_), .B(KEYINPUT36), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n534_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n578_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n583_), .A2(new_n577_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT71), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n580_), .A2(new_n584_), .A3(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n592_), .A3(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n534_), .A3(new_n591_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n600_), .A2(KEYINPUT72), .A3(new_n591_), .A4(new_n534_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n594_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G57gat), .B(G64gat), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(KEYINPUT11), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(KEYINPUT11), .ZN(new_n608_));
  XOR2_X1   g407(.A(G71gat), .B(G78gat), .Z(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n574_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n612_), .B(new_n550_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n574_), .A2(new_n613_), .A3(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .A4(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n614_), .A2(new_n618_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n617_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT5), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n629_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n621_), .A2(new_n624_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT13), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(KEYINPUT13), .A3(new_n632_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(G127gat), .B(G155gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT16), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G183gat), .B(G211gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(KEYINPUT73), .A2(KEYINPUT17), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT17), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(G231gat), .A2(G233gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n516_), .B(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(new_n612_), .ZN(new_n650_));
  MUX2_X1   g449(.A(new_n644_), .B(new_n647_), .S(new_n650_), .Z(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT74), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT74), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT75), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n605_), .A2(new_n638_), .A3(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n533_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n511_), .A3(new_n485_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n592_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n585_), .B2(KEYINPUT71), .ZN(new_n663_));
  AOI22_X1  g462(.A1(new_n663_), .A2(new_n599_), .B1(new_n590_), .B2(new_n586_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n505_), .A2(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n638_), .A2(new_n532_), .A3(new_n654_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G1gat), .B1(new_n667_), .B2(new_n445_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n659_), .A2(new_n660_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n661_), .A2(new_n668_), .A3(new_n669_), .ZN(G1324gat));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n665_), .A2(new_n323_), .A3(new_n666_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(new_n673_), .A3(G8gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n672_), .B2(G8gat), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT39), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n676_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n500_), .A2(G8gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n658_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n671_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n682_));
  AOI22_X1  g481(.A1(new_n675_), .A2(new_n676_), .B1(new_n658_), .B2(new_n679_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n675_), .A2(new_n676_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT40), .B(new_n683_), .C1(new_n684_), .C2(new_n674_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1325gat));
  OAI21_X1  g485(.A(G15gat), .B1(new_n667_), .B2(new_n455_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT41), .Z(new_n688_));
  INV_X1    g487(.A(G15gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n658_), .A2(new_n689_), .A3(new_n456_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1326gat));
  OAI21_X1  g490(.A(G22gat), .B1(new_n667_), .B2(new_n493_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT42), .ZN(new_n693_));
  INV_X1    g492(.A(G22gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n658_), .A2(new_n694_), .A3(new_n405_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1327gat));
  NAND2_X1  g495(.A1(new_n656_), .A2(new_n664_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(new_n638_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n533_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n445_), .A2(G29gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT109), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n603_), .A2(new_n604_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n594_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n505_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT102), .B1(new_n492_), .B2(new_n493_), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n459_), .B(new_n405_), .C1(new_n489_), .C2(new_n491_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n503_), .A2(new_n496_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n456_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n710_), .B(new_n605_), .C1(new_n715_), .C2(new_n458_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n709_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n637_), .A2(new_n531_), .A3(new_n656_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT106), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n717_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n722_), .B(new_n719_), .C1(new_n709_), .C2(new_n716_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n721_), .A2(new_n723_), .A3(new_n445_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G29gat), .B1(new_n724_), .B2(KEYINPUT107), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n721_), .A2(new_n723_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(KEYINPUT107), .A3(new_n485_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n705_), .B1(new_n725_), .B2(new_n727_), .ZN(G1328gat));
  INV_X1    g527(.A(G36gat), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n533_), .A2(new_n700_), .A3(new_n729_), .A4(new_n323_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT45), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n721_), .A2(new_n723_), .A3(new_n500_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT46), .B(new_n731_), .C1(new_n732_), .C2(new_n729_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n730_), .B(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n458_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n503_), .A2(new_n496_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n737_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n738_), .B2(new_n456_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n710_), .B1(new_n739_), .B2(new_n605_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n505_), .A2(new_n708_), .A3(KEYINPUT43), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n720_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n722_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n717_), .A2(KEYINPUT44), .A3(new_n720_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n323_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n735_), .B1(new_n745_), .B2(G36gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n733_), .B1(new_n746_), .B2(new_n747_), .ZN(G1329gat));
  NAND4_X1  g547(.A1(new_n743_), .A2(G43gat), .A3(new_n456_), .A4(new_n744_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n452_), .B1(new_n701_), .B2(new_n455_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(KEYINPUT47), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT47), .B1(new_n749_), .B2(new_n750_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1330gat));
  AOI21_X1  g552(.A(G50gat), .B1(new_n702_), .B2(new_n405_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n405_), .A2(G50gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n726_), .B2(new_n755_), .ZN(G1331gat));
  NOR3_X1   g555(.A1(new_n605_), .A2(new_n637_), .A3(new_n656_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(KEYINPUT111), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT111), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n505_), .A2(new_n531_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G57gat), .B1(new_n762_), .B2(new_n485_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n637_), .A2(new_n656_), .A3(new_n531_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n665_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(G57gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n485_), .B2(KEYINPUT112), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(KEYINPUT112), .B2(new_n766_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n763_), .B1(new_n765_), .B2(new_n768_), .ZN(G1332gat));
  NAND3_X1  g568(.A1(new_n665_), .A2(new_n323_), .A3(new_n764_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(G64gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G64gat), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n500_), .A2(G64gat), .ZN(new_n774_));
  OAI22_X1  g573(.A1(new_n772_), .A2(new_n773_), .B1(new_n761_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(G1333gat));
  INV_X1    g576(.A(G71gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n765_), .B2(new_n456_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT49), .Z(new_n780_));
  NAND3_X1  g579(.A1(new_n762_), .A2(new_n778_), .A3(new_n456_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1334gat));
  INV_X1    g581(.A(G78gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n765_), .B2(new_n405_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n785_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n405_), .A2(new_n783_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT115), .ZN(new_n789_));
  OAI22_X1  g588(.A1(new_n786_), .A2(new_n787_), .B1(new_n761_), .B2(new_n789_), .ZN(G1335gat));
  NAND3_X1  g589(.A1(new_n638_), .A2(new_n532_), .A3(new_n656_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n709_), .B2(new_n716_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793_), .B2(new_n445_), .ZN(new_n794_));
  NOR4_X1   g593(.A1(new_n505_), .A2(new_n699_), .A3(new_n531_), .A4(new_n637_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n544_), .A3(new_n485_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n793_), .B2(new_n500_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n545_), .A3(new_n323_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1337gat));
  INV_X1    g599(.A(new_n549_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n795_), .A2(new_n456_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n803_), .B(new_n535_), .C1(new_n792_), .C2(new_n456_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n791_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n456_), .B(new_n805_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT116), .B1(new_n806_), .B2(G99gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n802_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT51), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n802_), .C1(new_n804_), .C2(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1338gat));
  NAND3_X1  g611(.A1(new_n795_), .A2(new_n536_), .A3(new_n405_), .ZN(new_n813_));
  AOI211_X1 g612(.A(KEYINPUT52), .B(new_n536_), .C1(new_n792_), .C2(new_n405_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n405_), .B(new_n805_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(G106gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n814_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT53), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n813_), .C1(new_n814_), .C2(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1339gat));
  NOR3_X1   g621(.A1(new_n407_), .A2(new_n445_), .A3(new_n455_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(KEYINPUT59), .ZN(new_n825_));
  INV_X1    g624(.A(new_n656_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n621_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT55), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n621_), .A2(new_n827_), .A3(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n620_), .A2(new_n618_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n617_), .B1(new_n832_), .B2(new_n616_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n831_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n629_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT56), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n838_), .A3(new_n629_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n517_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n522_), .A2(new_n520_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n529_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n525_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n529_), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n844_), .B(KEYINPUT119), .Z(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n632_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n837_), .A2(KEYINPUT58), .A3(new_n839_), .A4(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n833_), .B1(new_n828_), .B2(KEYINPUT55), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n631_), .B1(new_n851_), .B2(new_n831_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n846_), .B1(new_n852_), .B2(new_n838_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n853_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n837_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n847_), .A2(new_n839_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n852_), .A2(new_n838_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n605_), .A2(new_n850_), .A3(new_n854_), .A4(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n632_), .A2(new_n531_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(KEYINPUT56), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n852_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n863_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n836_), .A2(new_n865_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n864_), .A2(new_n866_), .B1(new_n633_), .B2(new_n845_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n860_), .B1(new_n867_), .B2(new_n664_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n859_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n864_), .A2(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n633_), .A2(new_n845_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n664_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(KEYINPUT57), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT121), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n664_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(KEYINPUT57), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n826_), .B1(new_n869_), .B2(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n708_), .A2(new_n532_), .A3(new_n637_), .A4(new_n826_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT54), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n657_), .A2(new_n883_), .A3(new_n532_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n825_), .B1(new_n880_), .B2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n877_), .B1(new_n876_), .B2(KEYINPUT57), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n867_), .A2(KEYINPUT121), .A3(new_n860_), .A4(new_n664_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n859_), .A2(new_n868_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n654_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n882_), .A2(new_n884_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n824_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n886_), .B(new_n531_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(G113gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n891_), .A2(new_n892_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n823_), .ZN(new_n898_));
  OR3_X1    g697(.A1(new_n898_), .A2(G113gat), .A3(new_n532_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(G1340gat));
  OAI211_X1 g699(.A(new_n886_), .B(new_n638_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G120gat), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903_));
  AOI21_X1  g702(.A(G120gat), .B1(new_n638_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT122), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(KEYINPUT122), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n903_), .B2(G120gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n893_), .A2(new_n905_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n902_), .A2(new_n908_), .ZN(G1341gat));
  AOI21_X1  g708(.A(G127gat), .B1(new_n893_), .B2(new_n826_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n656_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n892_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n898_), .A2(KEYINPUT59), .B1(new_n912_), .B2(new_n825_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT123), .B(G127gat), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n654_), .A2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n910_), .B1(new_n913_), .B2(new_n915_), .ZN(G1342gat));
  OAI211_X1 g715(.A(new_n886_), .B(new_n605_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G134gat), .ZN(new_n918_));
  OR3_X1    g717(.A1(new_n898_), .A2(G134gat), .A3(new_n873_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1343gat));
  NOR4_X1   g719(.A1(new_n323_), .A2(new_n493_), .A3(new_n445_), .A4(new_n456_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n897_), .A2(new_n531_), .A3(new_n921_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g722(.A1(new_n897_), .A2(new_n638_), .A3(new_n921_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g724(.A1(new_n897_), .A2(new_n826_), .A3(new_n921_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT61), .B(G155gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1346gat));
  NAND2_X1  g727(.A1(new_n897_), .A2(new_n921_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G162gat), .B1(new_n929_), .B2(new_n708_), .ZN(new_n930_));
  OR2_X1    g729(.A1(new_n873_), .A2(G162gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(new_n931_), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n500_), .A2(new_n457_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n531_), .ZN(new_n934_));
  XOR2_X1   g733(.A(new_n934_), .B(KEYINPUT124), .Z(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n405_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n912_), .A2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n937_), .A2(new_n938_), .A3(G169gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n937_), .B2(G169gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n500_), .A2(new_n405_), .A3(new_n457_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n912_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n531_), .A2(new_n267_), .ZN(new_n943_));
  XOR2_X1   g742(.A(new_n943_), .B(KEYINPUT125), .Z(new_n944_));
  OAI22_X1  g743(.A1(new_n939_), .A2(new_n940_), .B1(new_n942_), .B2(new_n944_), .ZN(G1348gat));
  INV_X1    g744(.A(new_n942_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n638_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n869_), .A2(new_n879_), .ZN(new_n948_));
  AOI22_X1  g747(.A1(new_n948_), .A2(new_n654_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n405_), .ZN(new_n950_));
  AND3_X1   g749(.A1(new_n638_), .A2(G176gat), .A3(new_n933_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n947_), .A2(new_n266_), .B1(new_n950_), .B2(new_n951_), .ZN(G1349gat));
  AOI21_X1  g751(.A(new_n654_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n897_), .A2(new_n493_), .A3(new_n826_), .A4(new_n933_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n946_), .A2(new_n953_), .B1(new_n954_), .B2(new_n238_), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n942_), .B2(new_n708_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n664_), .A2(new_n241_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n942_), .B2(new_n957_), .ZN(G1351gat));
  NAND3_X1  g757(.A1(new_n502_), .A2(new_n323_), .A3(new_n455_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n949_), .A2(new_n959_), .ZN(new_n960_));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960_), .B2(new_n531_), .ZN(new_n961_));
  NOR4_X1   g760(.A1(new_n949_), .A2(new_n218_), .A3(new_n532_), .A4(new_n959_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1352gat));
  XNOR2_X1  g762(.A(KEYINPUT126), .B(G204gat), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n964_), .B1(new_n960_), .B2(new_n638_), .ZN(new_n965_));
  INV_X1    g764(.A(new_n964_), .ZN(new_n966_));
  NOR4_X1   g765(.A1(new_n949_), .A2(new_n637_), .A3(new_n959_), .A4(new_n966_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n965_), .A2(new_n967_), .ZN(G1353gat));
  NOR2_X1   g767(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(KEYINPUT127), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n654_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n970_), .B1(new_n960_), .B2(new_n971_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n970_), .ZN(new_n973_));
  INV_X1    g772(.A(new_n971_), .ZN(new_n974_));
  NOR4_X1   g773(.A1(new_n949_), .A2(new_n959_), .A3(new_n973_), .A4(new_n974_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n972_), .A2(new_n975_), .ZN(G1354gat));
  NAND3_X1  g775(.A1(new_n960_), .A2(new_n208_), .A3(new_n664_), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n949_), .A2(new_n708_), .A3(new_n959_), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n977_), .B1(new_n208_), .B2(new_n978_), .ZN(G1355gat));
endmodule


