//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n979_, new_n980_, new_n981_, new_n983_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n995_, new_n996_, new_n997_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1013_, new_n1014_, new_n1015_, new_n1017_, new_n1018_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1027_,
    new_n1028_, new_n1029_, new_n1031_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_;
  XNOR2_X1  g000(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n202_));
  AND2_X1   g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT75), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n205_), .B1(new_n207_), .B2(KEYINPUT78), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G106gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT64), .B1(new_n210_), .B2(new_n211_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n209_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G85gat), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT9), .A3(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n224_), .A2(KEYINPUT6), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(KEYINPUT6), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n216_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  INV_X1    g030(.A(G99gat), .ZN(new_n232_));
  INV_X1    g031(.A(G106gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n230_), .B(new_n234_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n219_), .A2(new_n220_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n236_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n229_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G43gat), .B(G50gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n245_), .A2(KEYINPUT15), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT15), .B1(new_n245_), .B2(new_n247_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n240_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n252_), .A2(new_n238_), .B1(new_n216_), .B2(new_n228_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n247_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n208_), .A2(new_n251_), .A3(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n207_), .A2(KEYINPUT78), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n259_), .A2(new_n208_), .A3(new_n251_), .A4(new_n255_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n261_), .A2(KEYINPUT79), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G190gat), .B(G218gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT76), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT77), .ZN(new_n265_));
  XOR2_X1   g064(.A(G134gat), .B(G162gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT36), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n268_), .B1(new_n261_), .B2(KEYINPUT79), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n267_), .A2(KEYINPUT36), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n262_), .A2(new_n269_), .B1(new_n270_), .B2(new_n261_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT104), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT24), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT24), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n278_), .B2(new_n274_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(new_n281_), .B2(G190gat), .ZN(new_n282_));
  INV_X1    g081(.A(G183gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT25), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G183gat), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n282_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G190gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT26), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n281_), .A2(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT84), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n279_), .B1(new_n287_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(G183gat), .A3(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT86), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT86), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n297_), .A2(new_n294_), .A3(G183gat), .A4(G190gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n299_), .A2(KEYINPUT85), .A3(KEYINPUT23), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT85), .B1(new_n299_), .B2(KEYINPUT23), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n296_), .B(new_n298_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n293_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G176gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT87), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT87), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G176gat), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT22), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT22), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G169gat), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n305_), .A2(new_n307_), .A3(new_n309_), .A4(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n312_), .A2(new_n277_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n299_), .A2(KEYINPUT23), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n295_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n303_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT30), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT88), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n322_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G71gat), .B(G99gat), .ZN(new_n325_));
  INV_X1    g124(.A(G43gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(G15gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n327_), .B(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n323_), .A2(new_n324_), .A3(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n324_), .A2(new_n330_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G127gat), .B(G134gat), .Z(new_n333_));
  XOR2_X1   g132(.A(G113gat), .B(G120gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT31), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n336_), .B(KEYINPUT89), .Z(new_n337_));
  NAND4_X1  g136(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT90), .A4(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT90), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n338_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G8gat), .B(G36gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT18), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT20), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n312_), .A2(new_n277_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(new_n317_), .B2(new_n302_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n289_), .A2(new_n290_), .A3(new_n284_), .A4(new_n286_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n274_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(KEYINPUT24), .A3(new_n277_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT100), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n352_), .A2(new_n354_), .A3(KEYINPUT100), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n315_), .A2(new_n276_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n351_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G218gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(G211gat), .ZN(new_n363_));
  INV_X1    g162(.A(G211gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G218gat), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n363_), .A2(new_n365_), .A3(KEYINPUT96), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT96), .B1(new_n363_), .B2(new_n365_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT21), .ZN(new_n369_));
  AND2_X1   g168(.A1(G197gat), .A2(G204gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(G197gat), .A2(G204gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G197gat), .ZN(new_n373_));
  INV_X1    g172(.A(G204gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G197gat), .A2(G204gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(KEYINPUT21), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n372_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n368_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT97), .B1(new_n370_), .B2(new_n371_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT97), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n375_), .A2(new_n381_), .A3(new_n376_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n380_), .A2(new_n382_), .A3(KEYINPUT21), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT98), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n368_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT96), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n364_), .A2(G218gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n362_), .A2(G211gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n363_), .A2(new_n365_), .A3(KEYINPUT96), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n380_), .A2(new_n382_), .A3(KEYINPUT21), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT98), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n379_), .B1(new_n385_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n349_), .B1(new_n361_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n385_), .A2(new_n393_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n379_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n320_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n395_), .A2(new_n398_), .A3(new_n402_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n293_), .A2(new_n302_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n349_), .B1(new_n394_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n358_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT100), .B1(new_n352_), .B2(new_n354_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n360_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n351_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n401_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n398_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n348_), .B1(new_n403_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n399_), .A2(new_n404_), .A3(new_n400_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT20), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n361_), .A2(new_n394_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n397_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n395_), .A2(new_n402_), .A3(new_n398_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n347_), .A3(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G85gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT0), .B(G57gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n335_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT91), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT92), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n434_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT2), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(G141gat), .B2(G148gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G141gat), .A2(G148gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(KEYINPUT2), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n439_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT93), .B1(new_n436_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(KEYINPUT2), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n440_), .A2(G141gat), .A3(G148gat), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n446_), .A2(new_n447_), .B1(new_n438_), .B2(new_n437_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n433_), .A2(new_n435_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT93), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n431_), .B1(new_n445_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n442_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(new_n437_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n429_), .B1(new_n428_), .B2(KEYINPUT1), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n426_), .B(KEYINPUT91), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT1), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n455_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n425_), .B1(new_n452_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n431_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n450_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n428_), .A2(KEYINPUT1), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n459_), .A2(new_n466_), .A3(new_n430_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n454_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n468_), .A3(new_n335_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G225gat), .A2(G233gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n461_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n461_), .A2(KEYINPUT4), .A3(new_n469_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n470_), .B1(new_n461_), .B2(KEYINPUT4), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n424_), .B(new_n472_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n413_), .A2(new_n419_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n461_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n471_), .B1(new_n461_), .B2(KEYINPUT4), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n477_), .B(new_n423_), .C1(new_n473_), .C2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT102), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n335_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT4), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n470_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n461_), .A2(KEYINPUT4), .A3(new_n469_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n487_), .A2(KEYINPUT102), .A3(new_n477_), .A4(new_n423_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n481_), .A2(new_n482_), .A3(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n424_), .A2(new_n482_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n487_), .A2(new_n477_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT101), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT101), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n487_), .A2(new_n493_), .A3(new_n477_), .A4(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n476_), .A2(new_n489_), .A3(new_n495_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n415_), .A2(new_n416_), .A3(new_n397_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n398_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n498_));
  OAI211_X1 g297(.A(KEYINPUT32), .B(new_n347_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n347_), .A2(KEYINPUT32), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n417_), .A2(new_n418_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n479_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n423_), .B1(new_n487_), .B2(new_n477_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n499_), .B(new_n501_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G22gat), .B(G50gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT29), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n465_), .A2(new_n468_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT28), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n465_), .A2(new_n468_), .A3(new_n509_), .A4(new_n506_), .ZN(new_n510_));
  INV_X1    g309(.A(G228gat), .ZN(new_n511_));
  INV_X1    g310(.A(G233gat), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n512_), .A2(KEYINPUT94), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(KEYINPUT94), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n511_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT95), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT99), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n508_), .A2(new_n510_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n505_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n445_), .A2(new_n451_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n460_), .B1(new_n523_), .B2(new_n462_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n509_), .B1(new_n524_), .B2(new_n506_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n510_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n518_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n505_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n508_), .A2(new_n510_), .A3(new_n519_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n516_), .A2(new_n517_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n401_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n506_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n533_));
  OAI21_X1  g332(.A(G78gat), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n399_), .A2(new_n400_), .B1(new_n517_), .B2(new_n516_), .ZN(new_n535_));
  INV_X1    g334(.A(G78gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT29), .B1(new_n452_), .B2(new_n460_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n534_), .A2(G106gat), .A3(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n536_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n233_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n522_), .A2(new_n530_), .A3(new_n539_), .A4(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n539_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n520_), .A2(new_n521_), .A3(new_n505_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n528_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n496_), .A2(new_n504_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(KEYINPUT103), .B(KEYINPUT27), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n417_), .A2(new_n347_), .A3(new_n418_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n347_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n348_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(KEYINPUT27), .A3(new_n419_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n547_), .A2(new_n553_), .A3(new_n543_), .A4(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n502_), .A2(new_n503_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n273_), .B(new_n343_), .C1(new_n548_), .C2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n553_), .A2(new_n555_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n547_), .A2(new_n543_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n343_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n557_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n560_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n561_), .A3(new_n557_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n504_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n413_), .A2(new_n419_), .A3(new_n475_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n571_), .B2(new_n489_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n568_), .B1(new_n572_), .B2(new_n563_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n273_), .B1(new_n573_), .B2(new_n343_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT105), .B(new_n272_), .C1(new_n567_), .C2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n343_), .B1(new_n548_), .B2(new_n559_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT104), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n566_), .A3(new_n560_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT105), .B1(new_n579_), .B2(new_n272_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT72), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT71), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT66), .B(G71gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(G78gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n536_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(G64gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(G57gat), .ZN(new_n590_));
  INV_X1    g389(.A(G57gat), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(G64gat), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n590_), .A2(new_n592_), .A3(KEYINPUT11), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT11), .B1(new_n590_), .B2(new_n592_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n585_), .B(new_n588_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(new_n592_), .A3(KEYINPUT11), .ZN(new_n596_));
  INV_X1    g395(.A(new_n588_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n536_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT67), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n595_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT68), .B1(new_n603_), .B2(new_n241_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(new_n599_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT67), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n595_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n241_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT68), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n253_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n608_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n608_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n614_), .B1(new_n609_), .B2(new_n253_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n605_), .A2(KEYINPUT69), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT69), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n241_), .B(KEYINPUT12), .C1(new_n619_), .C2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(G120gat), .B(G148gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n615_), .A2(new_n623_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n615_), .B2(new_n623_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n583_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n615_), .A2(new_n623_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n615_), .A2(new_n623_), .A3(new_n628_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(KEYINPUT71), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n582_), .B1(new_n637_), .B2(KEYINPUT13), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT13), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n631_), .A2(new_n636_), .A3(KEYINPUT72), .A4(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT73), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n637_), .B2(KEYINPUT13), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n637_), .A2(new_n642_), .A3(KEYINPUT13), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(G229gat), .A2(G233gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G1gat), .B(G8gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT81), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT80), .B(G1gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G8gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT14), .ZN(new_n653_));
  XOR2_X1   g452(.A(G15gat), .B(G22gat), .Z(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n650_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT14), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n651_), .B2(G8gat), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n658_), .A2(KEYINPUT81), .A3(new_n654_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n649_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n653_), .A2(new_n650_), .A3(new_n655_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT81), .B1(new_n658_), .B2(new_n654_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n648_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(new_n254_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n254_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n647_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n660_), .A2(new_n250_), .A3(new_n663_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT82), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT82), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n660_), .A2(new_n250_), .A3(new_n663_), .A4(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n669_), .A2(new_n666_), .A3(new_n647_), .A4(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT83), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n667_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(KEYINPUT83), .ZN(new_n676_));
  XNOR2_X1  g475(.A(G113gat), .B(G141gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(G169gat), .B(G197gat), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n677_), .B(new_n678_), .Z(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n676_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n679_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n647_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n666_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n664_), .A2(new_n254_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(new_n672_), .B2(KEYINPUT83), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n672_), .A2(KEYINPUT83), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n681_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n680_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n646_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n664_), .ZN(new_n691_));
  AND2_X1   g490(.A1(G231gat), .A2(G233gat), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n692_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n619_), .A2(new_n621_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n696_), .ZN(new_n698_));
  XOR2_X1   g497(.A(G127gat), .B(G155gat), .Z(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT16), .ZN(new_n700_));
  XNOR2_X1  g499(.A(G183gat), .B(G211gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT17), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n697_), .A2(new_n698_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n695_), .A2(new_n609_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n693_), .A2(new_n603_), .A3(new_n694_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n702_), .B(KEYINPUT17), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n690_), .A2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n581_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n558_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G1gat), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n579_), .A2(new_n689_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n710_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n261_), .A2(new_n270_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n717_), .B(KEYINPUT37), .C1(new_n261_), .C2(new_n268_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n716_), .B(new_n718_), .C1(new_n271_), .C2(KEYINPUT37), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n637_), .A2(KEYINPUT13), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT73), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n644_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n719_), .B1(new_n722_), .B2(new_n641_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n715_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n651_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n558_), .A3(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT38), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n714_), .A2(new_n727_), .ZN(G1324gat));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n562_), .B(new_n711_), .C1(new_n576_), .C2(new_n580_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(G8gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n730_), .B2(G8gat), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT39), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n730_), .A2(G8gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(KEYINPUT106), .A3(new_n734_), .ZN(new_n737_));
  INV_X1    g536(.A(G8gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n724_), .A2(new_n738_), .A3(new_n562_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n729_), .B1(new_n735_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(KEYINPUT106), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n730_), .A2(new_n731_), .A3(G8gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(KEYINPUT39), .A3(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n744_), .A2(KEYINPUT40), .A3(new_n737_), .A4(new_n739_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n741_), .A2(new_n745_), .ZN(G1325gat));
  NAND2_X1  g545(.A1(new_n712_), .A2(new_n565_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G15gat), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT41), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT41), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(new_n750_), .A3(G15gat), .ZN(new_n751_));
  INV_X1    g550(.A(G15gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n724_), .A2(new_n752_), .A3(new_n565_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT107), .Z(new_n754_));
  NAND3_X1  g553(.A1(new_n749_), .A2(new_n751_), .A3(new_n754_), .ZN(G1326gat));
  INV_X1    g554(.A(G22gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n724_), .A2(new_n756_), .A3(new_n563_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n712_), .A2(new_n563_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(G22gat), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT42), .B(new_n756_), .C1(new_n712_), .C2(new_n563_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1327gat));
  AOI22_X1  g561(.A1(new_n721_), .A2(new_n644_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n271_), .A2(new_n710_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n715_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G29gat), .B1(new_n766_), .B2(new_n558_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n646_), .A2(new_n689_), .A3(new_n710_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n718_), .B1(new_n271_), .B2(KEYINPUT37), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n770_), .B(new_n771_), .C1(new_n567_), .C2(new_n574_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n770_), .B1(new_n579_), .B2(new_n771_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n769_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT108), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n771_), .B1(new_n567_), .B2(new_n574_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT43), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n772_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n769_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n777_), .A3(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n769_), .B(KEYINPUT44), .C1(new_n773_), .C2(new_n774_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n558_), .A2(G29gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n767_), .B1(new_n785_), .B2(new_n786_), .ZN(G1328gat));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT46), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT110), .Z(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(G36gat), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n784_), .A2(new_n562_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n783_), .B2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n788_), .A2(KEYINPUT46), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n561_), .A2(G36gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n766_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n715_), .A2(new_n765_), .A3(new_n798_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT45), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n796_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n791_), .B1(new_n795_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT44), .B1(new_n775_), .B2(KEYINPUT108), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n793_), .B1(new_n805_), .B2(new_n782_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n790_), .B(new_n802_), .C1(new_n806_), .C2(new_n792_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(G1329gat));
  NAND2_X1  g607(.A1(new_n565_), .A2(G43gat), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n768_), .B1(new_n779_), .B2(new_n772_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n777_), .B1(new_n811_), .B2(new_n781_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n775_), .A2(KEYINPUT108), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n784_), .B(new_n810_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n715_), .A2(new_n565_), .A3(new_n765_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n326_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n815_), .B2(new_n326_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n814_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT47), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n814_), .A2(new_n822_), .A3(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1330gat));
  AOI21_X1  g623(.A(G50gat), .B1(new_n766_), .B2(new_n563_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n563_), .A2(G50gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n785_), .B2(new_n826_), .ZN(G1331gat));
  NOR3_X1   g626(.A1(new_n646_), .A2(new_n689_), .A3(new_n710_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n581_), .A2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n557_), .A2(new_n591_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n689_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n579_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n719_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n763_), .A2(new_n834_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT112), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n557_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G57gat), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT113), .B1(new_n831_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n838_), .A2(new_n840_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n843_), .A2(new_n591_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(G1332gat));
  NAND3_X1  g646(.A1(new_n837_), .A2(new_n589_), .A3(new_n562_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT48), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n829_), .A2(new_n562_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(G64gat), .ZN(new_n851_));
  AOI211_X1 g650(.A(KEYINPUT48), .B(new_n589_), .C1(new_n829_), .C2(new_n562_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n848_), .B1(new_n851_), .B2(new_n852_), .ZN(G1333gat));
  OR3_X1    g652(.A1(new_n836_), .A2(G71gat), .A3(new_n343_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n829_), .A2(new_n565_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n855_), .A2(G71gat), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n855_), .B2(G71gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n857_), .B2(new_n858_), .ZN(G1334gat));
  NAND3_X1  g658(.A1(new_n837_), .A2(new_n536_), .A3(new_n563_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n829_), .A2(new_n563_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(G78gat), .ZN(new_n863_));
  AOI211_X1 g662(.A(KEYINPUT50), .B(new_n536_), .C1(new_n829_), .C2(new_n563_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n860_), .B1(new_n863_), .B2(new_n864_), .ZN(G1335gat));
  NOR3_X1   g664(.A1(new_n833_), .A2(new_n646_), .A3(new_n764_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n217_), .A3(new_n558_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n716_), .A2(new_n689_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n763_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT115), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n763_), .A2(new_n871_), .A3(new_n868_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n780_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n558_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n867_), .B1(new_n876_), .B2(new_n217_), .ZN(G1336gat));
  NAND3_X1  g676(.A1(new_n866_), .A2(new_n218_), .A3(new_n562_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n562_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n880_), .B2(new_n218_), .ZN(G1337gat));
  AOI21_X1  g680(.A(new_n232_), .B1(new_n874_), .B2(new_n565_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n214_), .A2(new_n215_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n866_), .A2(new_n565_), .A3(new_n883_), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n882_), .A2(KEYINPUT51), .A3(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT51), .B1(new_n882_), .B2(new_n884_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1338gat));
  NAND3_X1  g686(.A1(new_n866_), .A2(new_n563_), .A3(new_n209_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n873_), .B(new_n563_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n889_), .A2(new_n890_), .A3(G106gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n889_), .B2(G106gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n888_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g693(.A1(new_n646_), .A2(new_n834_), .A3(new_n832_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT54), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n723_), .A2(new_n897_), .A3(new_n832_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n623_), .A2(KEYINPUT116), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT55), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT55), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n623_), .A2(KEYINPUT116), .A3(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n617_), .A2(new_n604_), .A3(new_n611_), .A4(new_n622_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n614_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n901_), .A2(new_n903_), .A3(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n633_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n906_), .A2(KEYINPUT56), .A3(new_n633_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n679_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n686_), .A2(new_n687_), .A3(new_n681_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n635_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n682_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n916_));
  OAI21_X1  g715(.A(KEYINPUT117), .B1(new_n916_), .B2(new_n679_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n669_), .A2(new_n666_), .A3(new_n682_), .A4(new_n671_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n647_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n919_), .A2(new_n920_), .A3(new_n681_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n917_), .A2(new_n918_), .A3(new_n921_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n680_), .A2(new_n922_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n911_), .A2(new_n915_), .B1(new_n637_), .B2(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n899_), .B1(new_n924_), .B2(new_n271_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n680_), .A2(new_n635_), .A3(new_n922_), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n906_), .A2(KEYINPUT56), .A3(new_n633_), .ZN(new_n927_));
  AOI21_X1  g726(.A(KEYINPUT56), .B1(new_n906_), .B2(new_n633_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT58), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n911_), .A2(KEYINPUT58), .A3(new_n926_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n931_), .A2(new_n932_), .A3(new_n771_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n899_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n914_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n637_), .A2(new_n923_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n272_), .B(new_n934_), .C1(new_n935_), .C2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n925_), .A2(new_n933_), .A3(new_n937_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n896_), .A2(new_n898_), .B1(new_n938_), .B2(new_n710_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n564_), .A2(new_n558_), .A3(new_n565_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(G113gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n941_), .A2(new_n942_), .A3(new_n689_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n944_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n933_), .A2(new_n937_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n911_), .A2(new_n915_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n637_), .A2(new_n923_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n934_), .B1(new_n949_), .B2(new_n272_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n710_), .B1(new_n946_), .B2(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n897_), .B1(new_n723_), .B2(new_n832_), .ZN(new_n952_));
  NOR4_X1   g751(.A1(new_n763_), .A2(KEYINPUT54), .A3(new_n689_), .A4(new_n719_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n951_), .B1(new_n952_), .B2(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n940_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n954_), .A2(KEYINPUT59), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n832_), .B1(new_n945_), .B2(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n943_), .B1(new_n957_), .B2(new_n942_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(KEYINPUT119), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n960_), .B(new_n943_), .C1(new_n957_), .C2(new_n942_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n959_), .A2(new_n961_), .ZN(G1340gat));
  INV_X1    g761(.A(G120gat), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n963_), .B1(new_n646_), .B2(KEYINPUT60), .ZN(new_n964_));
  OAI211_X1 g763(.A(new_n941_), .B(new_n964_), .C1(KEYINPUT60), .C2(new_n963_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(KEYINPUT120), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n945_), .A2(new_n956_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G120gat), .B1(new_n967_), .B2(new_n646_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n966_), .A2(new_n968_), .ZN(G1341gat));
  OAI21_X1  g768(.A(G127gat), .B1(new_n967_), .B2(new_n710_), .ZN(new_n970_));
  INV_X1    g769(.A(G127gat), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n941_), .A2(new_n971_), .A3(new_n716_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n970_), .A2(new_n972_), .ZN(G1342gat));
  INV_X1    g772(.A(new_n771_), .ZN(new_n974_));
  OAI21_X1  g773(.A(G134gat), .B1(new_n967_), .B2(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(G134gat), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n941_), .A2(new_n976_), .A3(new_n271_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n977_), .ZN(G1343gat));
  NOR3_X1   g777(.A1(new_n565_), .A2(new_n557_), .A3(new_n556_), .ZN(new_n979_));
  AND2_X1   g778(.A1(new_n954_), .A2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n980_), .A2(new_n689_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g781(.A1(new_n980_), .A2(new_n763_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(new_n983_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g783(.A1(new_n980_), .A2(new_n716_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n985_), .A2(KEYINPUT121), .ZN(new_n986_));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n987_));
  NAND3_X1  g786(.A1(new_n980_), .A2(new_n987_), .A3(new_n716_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n986_), .A2(new_n988_), .ZN(new_n989_));
  XNOR2_X1  g788(.A(KEYINPUT61), .B(G155gat), .ZN(new_n990_));
  INV_X1    g789(.A(new_n990_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n989_), .A2(new_n991_), .ZN(new_n992_));
  NAND3_X1  g791(.A1(new_n986_), .A2(new_n988_), .A3(new_n990_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n992_), .A2(new_n993_), .ZN(G1346gat));
  INV_X1    g793(.A(new_n980_), .ZN(new_n995_));
  OAI21_X1  g794(.A(G162gat), .B1(new_n995_), .B2(new_n974_), .ZN(new_n996_));
  OR2_X1    g795(.A1(new_n272_), .A2(G162gat), .ZN(new_n997_));
  OAI21_X1  g796(.A(new_n996_), .B1(new_n995_), .B2(new_n997_), .ZN(G1347gat));
  NOR4_X1   g797(.A1(new_n343_), .A2(new_n563_), .A3(new_n561_), .A4(new_n558_), .ZN(new_n999_));
  AND2_X1   g798(.A1(new_n954_), .A2(new_n999_), .ZN(new_n1000_));
  NAND3_X1  g799(.A1(new_n689_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n1001_));
  XOR2_X1   g800(.A(new_n1001_), .B(KEYINPUT123), .Z(new_n1002_));
  NAND2_X1  g801(.A1(new_n1000_), .A2(new_n1002_), .ZN(new_n1003_));
  NAND3_X1  g802(.A1(new_n954_), .A2(new_n689_), .A3(new_n999_), .ZN(new_n1004_));
  XOR2_X1   g803(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n1005_));
  AND3_X1   g804(.A1(new_n1004_), .A2(G169gat), .A3(new_n1005_), .ZN(new_n1006_));
  AOI21_X1  g805(.A(new_n1005_), .B1(new_n1004_), .B2(G169gat), .ZN(new_n1007_));
  OAI21_X1  g806(.A(new_n1003_), .B1(new_n1006_), .B2(new_n1007_), .ZN(new_n1008_));
  INV_X1    g807(.A(KEYINPUT124), .ZN(new_n1009_));
  NAND2_X1  g808(.A1(new_n1008_), .A2(new_n1009_), .ZN(new_n1010_));
  OAI211_X1 g809(.A(KEYINPUT124), .B(new_n1003_), .C1(new_n1006_), .C2(new_n1007_), .ZN(new_n1011_));
  NAND2_X1  g810(.A1(new_n1010_), .A2(new_n1011_), .ZN(G1348gat));
  NAND2_X1  g811(.A1(new_n1000_), .A2(new_n763_), .ZN(new_n1013_));
  NOR2_X1   g812(.A1(new_n1013_), .A2(new_n304_), .ZN(new_n1014_));
  AND2_X1   g813(.A1(new_n305_), .A2(new_n307_), .ZN(new_n1015_));
  AOI21_X1  g814(.A(new_n1014_), .B1(new_n1015_), .B2(new_n1013_), .ZN(G1349gat));
  NAND2_X1  g815(.A1(new_n1000_), .A2(new_n716_), .ZN(new_n1017_));
  AOI21_X1  g816(.A(new_n1017_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n1018_));
  AOI21_X1  g817(.A(new_n1018_), .B1(new_n283_), .B2(new_n1017_), .ZN(G1350gat));
  NOR2_X1   g818(.A1(new_n272_), .A2(new_n291_), .ZN(new_n1020_));
  AND2_X1   g819(.A1(new_n1000_), .A2(new_n1020_), .ZN(new_n1021_));
  AOI21_X1  g820(.A(new_n288_), .B1(new_n1000_), .B2(new_n771_), .ZN(new_n1022_));
  INV_X1    g821(.A(KEYINPUT125), .ZN(new_n1023_));
  OR3_X1    g822(.A1(new_n1021_), .A2(new_n1022_), .A3(new_n1023_), .ZN(new_n1024_));
  OAI21_X1  g823(.A(new_n1023_), .B1(new_n1021_), .B2(new_n1022_), .ZN(new_n1025_));
  NAND2_X1  g824(.A1(new_n1024_), .A2(new_n1025_), .ZN(G1351gat));
  NOR2_X1   g825(.A1(new_n565_), .A2(new_n558_), .ZN(new_n1027_));
  AND4_X1   g826(.A1(new_n563_), .A2(new_n954_), .A3(new_n562_), .A4(new_n1027_), .ZN(new_n1028_));
  NAND2_X1  g827(.A1(new_n1028_), .A2(new_n689_), .ZN(new_n1029_));
  XNOR2_X1  g828(.A(new_n1029_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g829(.A1(new_n1028_), .A2(new_n763_), .ZN(new_n1031_));
  XNOR2_X1  g830(.A(new_n1031_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g831(.A1(new_n1028_), .A2(new_n716_), .ZN(new_n1033_));
  XNOR2_X1  g832(.A(KEYINPUT63), .B(G211gat), .ZN(new_n1034_));
  NOR2_X1   g833(.A1(new_n1033_), .A2(new_n1034_), .ZN(new_n1035_));
  NOR2_X1   g834(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1036_));
  AOI21_X1  g835(.A(new_n1035_), .B1(new_n1033_), .B2(new_n1036_), .ZN(G1354gat));
  INV_X1    g836(.A(KEYINPUT126), .ZN(new_n1038_));
  NOR2_X1   g837(.A1(new_n272_), .A2(G218gat), .ZN(new_n1039_));
  NAND2_X1  g838(.A1(new_n1028_), .A2(new_n1039_), .ZN(new_n1040_));
  AND2_X1   g839(.A1(new_n1028_), .A2(new_n771_), .ZN(new_n1041_));
  OAI211_X1 g840(.A(new_n1038_), .B(new_n1040_), .C1(new_n1041_), .C2(new_n362_), .ZN(new_n1042_));
  INV_X1    g841(.A(new_n1040_), .ZN(new_n1043_));
  AOI21_X1  g842(.A(new_n362_), .B1(new_n1028_), .B2(new_n771_), .ZN(new_n1044_));
  OAI21_X1  g843(.A(KEYINPUT126), .B1(new_n1043_), .B2(new_n1044_), .ZN(new_n1045_));
  NAND2_X1  g844(.A1(new_n1042_), .A2(new_n1045_), .ZN(G1355gat));
endmodule


