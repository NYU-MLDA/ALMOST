//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n602_, new_n603_, new_n604_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT31), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT84), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n205_), .A2(new_n206_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(KEYINPUT84), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n204_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G227gat), .A2(G233gat), .ZN(new_n214_));
  INV_X1    g013(.A(G15gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT30), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n213_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT82), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n223_));
  OR3_X1    g022(.A1(new_n222_), .A2(new_n223_), .A3(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT23), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT23), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n220_), .B(new_n224_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT81), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(KEYINPUT24), .A3(new_n220_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n226_), .A2(KEYINPUT26), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT80), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n225_), .A2(KEYINPUT79), .A3(KEYINPUT25), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n226_), .A2(KEYINPUT26), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT25), .B1(new_n225_), .B2(KEYINPUT79), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n235_), .B1(new_n237_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n229_), .A2(KEYINPUT83), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT83), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n228_), .A2(new_n244_), .A3(KEYINPUT23), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n227_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(KEYINPUT24), .B2(new_n234_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n232_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT85), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n218_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n218_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G228gat), .A2(G233gat), .ZN(new_n255_));
  INV_X1    g054(.A(G78gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G106gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n260_), .A2(KEYINPUT1), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(KEYINPUT1), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(G141gat), .ZN(new_n266_));
  INV_X1    g065(.A(G148gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n264_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT87), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n266_), .A2(new_n267_), .A3(KEYINPUT3), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(G141gat), .B2(G148gat), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT2), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n276_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT86), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n272_), .A2(new_n274_), .ZN(new_n281_));
  AND3_X1   g080(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n260_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(new_n263_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n271_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  AOI211_X1 g090(.A(KEYINPUT87), .B(new_n291_), .C1(new_n280_), .C2(new_n286_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n270_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT28), .B1(new_n293_), .B2(KEYINPUT29), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT88), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n281_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n285_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n289_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT87), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n271_), .B(new_n289_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n269_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n294_), .A2(new_n295_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n295_), .B1(new_n294_), .B2(new_n304_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n259_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n259_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n305_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G211gat), .B(G218gat), .Z(new_n313_));
  INV_X1    g112(.A(G197gat), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT90), .ZN(new_n315_));
  INV_X1    g114(.A(G204gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(KEYINPUT90), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT21), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(G197gat), .B2(G204gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n313_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(G204gat), .A3(new_n317_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n316_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT91), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n314_), .B2(G204gat), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .A4(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n322_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n313_), .A2(KEYINPUT21), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT89), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT89), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n335_), .B(new_n332_), .C1(new_n301_), .C2(new_n303_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G22gat), .B(G50gat), .Z(new_n338_));
  OR2_X1    g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n338_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n312_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n339_), .A2(new_n308_), .A3(new_n311_), .A4(new_n340_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n207_), .A2(new_n209_), .ZN(new_n345_));
  AOI211_X1 g144(.A(new_n269_), .B(new_n345_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n212_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT95), .B1(new_n293_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT95), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n301_), .A2(new_n350_), .A3(new_n212_), .ZN(new_n351_));
  OAI211_X1 g150(.A(KEYINPUT4), .B(new_n347_), .C1(new_n349_), .C2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT96), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n350_), .B1(new_n301_), .B2(new_n212_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n293_), .A2(KEYINPUT95), .A3(new_n348_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n346_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT96), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(KEYINPUT4), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n301_), .A2(KEYINPUT4), .A3(new_n212_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n353_), .A2(new_n355_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n357_), .ZN(new_n363_));
  AND4_X1   g162(.A1(KEYINPUT97), .A2(new_n363_), .A3(new_n354_), .A4(new_n347_), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT97), .B1(new_n358_), .B2(new_n354_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G85gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT0), .B(G57gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  NAND3_X1  g169(.A1(new_n362_), .A2(new_n366_), .A3(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(KEYINPUT98), .B(KEYINPUT33), .Z(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n362_), .A2(new_n366_), .A3(KEYINPUT33), .A4(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT19), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n249_), .A2(new_n332_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT20), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n234_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT24), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n227_), .A2(new_n229_), .B1(new_n381_), .B2(new_n233_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n239_), .A2(new_n236_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT93), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT25), .B(G183gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n380_), .B(new_n382_), .C1(new_n384_), .C2(new_n386_), .ZN(new_n387_));
  OR3_X1    g186(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT94), .ZN(new_n388_));
  INV_X1    g187(.A(G176gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT94), .B1(new_n222_), .B2(new_n223_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n247_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n391_), .B(new_n220_), .C1(new_n392_), .C2(new_n231_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n387_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(new_n332_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n377_), .B1(new_n379_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n332_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n328_), .A2(new_n331_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n398_), .B(new_n232_), .C1(new_n248_), .C2(new_n242_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n397_), .A2(new_n399_), .A3(KEYINPUT20), .A4(new_n376_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT18), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n401_), .B(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n353_), .A2(new_n354_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n370_), .B1(new_n358_), .B2(new_n355_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n373_), .A2(new_n374_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT99), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n332_), .B1(new_n394_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n412_), .B2(new_n394_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n378_), .A2(KEYINPUT20), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n377_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AND4_X1   g215(.A1(KEYINPUT20), .A2(new_n397_), .A3(new_n377_), .A4(new_n399_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n401_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n406_), .A2(KEYINPUT32), .ZN(new_n420_));
  MUX2_X1   g219(.A(new_n418_), .B(new_n419_), .S(new_n420_), .Z(new_n421_));
  AND3_X1   g220(.A1(new_n362_), .A2(new_n366_), .A3(new_n370_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n370_), .B1(new_n362_), .B2(new_n366_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n344_), .B1(new_n411_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT100), .B1(new_n401_), .B2(new_n406_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT100), .ZN(new_n428_));
  AOI211_X1 g227(.A(new_n428_), .B(new_n405_), .C1(new_n396_), .C2(new_n400_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n405_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n426_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n407_), .A2(KEYINPUT27), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n342_), .B(new_n343_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n423_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n371_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n254_), .B1(new_n425_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n436_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n344_), .A2(new_n254_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n432_), .A2(new_n433_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G230gat), .A2(G233gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n444_), .B(KEYINPUT64), .Z(new_n445_));
  XNOR2_X1  g244(.A(G85gat), .B(G92gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT65), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(KEYINPUT8), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G99gat), .A2(G106gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n448_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT8), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(KEYINPUT65), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G85gat), .ZN(new_n458_));
  INV_X1    g257(.A(G92gat), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n458_), .A2(new_n459_), .A3(KEYINPUT9), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n451_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT9), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT10), .B(G99gat), .ZN(new_n463_));
  OAI221_X1 g262(.A(new_n461_), .B1(new_n462_), .B2(new_n446_), .C1(G106gat), .C2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n457_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n455_), .B1(KEYINPUT65), .B2(new_n456_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G57gat), .B(G64gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT11), .ZN(new_n469_));
  XOR2_X1   g268(.A(G71gat), .B(G78gat), .Z(new_n470_));
  OR2_X1    g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n468_), .A2(KEYINPUT11), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n470_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n467_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n467_), .A2(new_n474_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n445_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT66), .ZN(new_n479_));
  AND2_X1   g278(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n477_), .B1(new_n482_), .B2(new_n480_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n445_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT68), .B1(new_n475_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  AOI211_X1 g285(.A(new_n486_), .B(new_n445_), .C1(new_n467_), .C2(new_n474_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n481_), .B(new_n483_), .C1(new_n485_), .C2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n479_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G120gat), .B(G148gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT5), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n493_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n479_), .A2(new_n488_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT13), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(KEYINPUT13), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n497_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n501_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G1gat), .B(G8gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT74), .ZN(new_n507_));
  INV_X1    g306(.A(G22gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n215_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G15gat), .A2(G22gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G1gat), .A2(G8gat), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n509_), .A2(new_n510_), .B1(KEYINPUT14), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n507_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G29gat), .B(G36gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT77), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n513_), .A2(new_n516_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n507_), .B(new_n512_), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n516_), .B(KEYINPUT15), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n513_), .A2(new_n516_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n520_), .A3(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n527_), .A2(KEYINPUT78), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(KEYINPUT78), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n522_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n522_), .A2(new_n528_), .A3(new_n529_), .A4(new_n533_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n505_), .A2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n443_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G190gat), .B(G218gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT70), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n545_), .A2(KEYINPUT36), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT71), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT72), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n467_), .A2(new_n516_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n524_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n549_), .B(new_n550_), .C1(KEYINPUT35), .C2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n544_), .B(KEYINPUT36), .Z(new_n557_));
  OR2_X1    g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n559_), .A2(KEYINPUT37), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n557_), .B(KEYINPUT73), .Z(new_n561_));
  OAI21_X1  g360(.A(new_n556_), .B1(new_n555_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT37), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n474_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n523_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT75), .ZN(new_n569_));
  XOR2_X1   g368(.A(G127gat), .B(G155gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT16), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT17), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT76), .Z(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n568_), .A2(new_n577_), .A3(new_n573_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n565_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n540_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(G1gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n436_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT38), .ZN(new_n584_));
  INV_X1    g383(.A(new_n559_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n540_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(G1gat), .B1(new_n587_), .B2(new_n439_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(G1324gat));
  OAI21_X1  g388(.A(G8gat), .B1(new_n587_), .B2(new_n441_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT101), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT39), .B1(new_n590_), .B2(new_n591_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G8gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n441_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n581_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n592_), .A2(new_n593_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g400(.A(G15gat), .B1(new_n587_), .B2(new_n254_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT41), .Z(new_n603_));
  NAND3_X1  g402(.A1(new_n581_), .A2(new_n215_), .A3(new_n253_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(G1326gat));
  INV_X1    g404(.A(new_n344_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G22gat), .B1(new_n587_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n581_), .A2(new_n508_), .A3(new_n344_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1327gat));
  INV_X1    g410(.A(new_n579_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(new_n559_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n540_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(G29gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n436_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT44), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(KEYINPUT103), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT43), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n443_), .B2(new_n565_), .ZN(new_n621_));
  AOI211_X1 g420(.A(KEYINPUT43), .B(new_n564_), .C1(new_n438_), .C2(new_n442_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n612_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n539_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n619_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n619_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n627_), .B(new_n628_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n439_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n616_), .B1(new_n630_), .B2(new_n615_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT105), .Z(G1328gat));
  INV_X1    g431(.A(G36gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n614_), .A2(new_n633_), .A3(new_n596_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT45), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n443_), .A2(new_n565_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT43), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n443_), .A2(new_n620_), .A3(new_n565_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n628_), .B1(new_n640_), .B2(new_n627_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n629_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n636_), .B(new_n596_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G36gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n626_), .A2(new_n629_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n636_), .B1(new_n645_), .B2(new_n596_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n635_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT107), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(KEYINPUT107), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n645_), .A2(new_n596_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT106), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n441_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n633_), .B1(new_n654_), .B2(new_n636_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n656_), .A2(KEYINPUT107), .A3(new_n648_), .A4(new_n635_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n651_), .A2(new_n657_), .ZN(G1329gat));
  AOI21_X1  g457(.A(G43gat), .B1(new_n614_), .B2(new_n253_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n253_), .A2(G43gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n645_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(G1330gat));
  INV_X1    g462(.A(G50gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n344_), .A2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT110), .Z(new_n666_));
  NAND2_X1  g465(.A1(new_n614_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n645_), .A2(new_n344_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(G50gat), .ZN(new_n670_));
  AOI211_X1 g469(.A(KEYINPUT109), .B(new_n664_), .C1(new_n645_), .C2(new_n344_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT111), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT111), .B(new_n667_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1331gat));
  INV_X1    g475(.A(new_n505_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n537_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(new_n443_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n580_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT112), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT112), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n436_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(G57gat), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n679_), .A2(new_n586_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n439_), .A2(new_n685_), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n684_), .A2(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(G1332gat));
  INV_X1    g487(.A(G64gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n686_), .B2(new_n596_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n681_), .A2(new_n689_), .A3(new_n596_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1333gat));
  INV_X1    g493(.A(G71gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n686_), .B2(new_n253_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n681_), .A2(new_n695_), .A3(new_n253_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1334gat));
  AOI21_X1  g499(.A(new_n256_), .B1(new_n686_), .B2(new_n344_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT50), .Z(new_n702_));
  NAND3_X1  g501(.A1(new_n681_), .A2(new_n256_), .A3(new_n344_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1335gat));
  AND2_X1   g503(.A1(new_n679_), .A2(new_n613_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n458_), .A3(new_n436_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n640_), .A2(new_n579_), .A3(new_n678_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n436_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n710_), .B2(new_n458_), .ZN(G1336gat));
  OAI21_X1  g510(.A(G92gat), .B1(new_n707_), .B2(new_n441_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n705_), .A2(new_n459_), .A3(new_n596_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT115), .Z(G1337gat));
  OAI21_X1  g514(.A(G99gat), .B1(new_n707_), .B2(new_n254_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n463_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n705_), .A2(new_n717_), .A3(new_n253_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n719_), .B(new_n720_), .Z(G1338gat));
  AOI21_X1  g520(.A(new_n258_), .B1(new_n708_), .B2(new_n344_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n722_), .A2(KEYINPUT52), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(KEYINPUT52), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n705_), .A2(new_n258_), .A3(new_n344_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT117), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(new_n724_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT53), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT53), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n723_), .A2(new_n729_), .A3(new_n724_), .A4(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1339gat));
  INV_X1    g530(.A(KEYINPUT121), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT58), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n519_), .A2(new_n520_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n525_), .A2(new_n521_), .A3(new_n526_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n534_), .A3(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n536_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n496_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT120), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n485_), .A2(new_n487_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n740_), .A2(KEYINPUT55), .A3(new_n483_), .A4(new_n481_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n488_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n481_), .A2(new_n483_), .A3(new_n475_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n445_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n741_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(KEYINPUT56), .A3(new_n493_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT56), .B1(new_n746_), .B2(new_n493_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n733_), .B1(new_n739_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n565_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n739_), .A2(new_n733_), .A3(new_n750_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n749_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT118), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n747_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n749_), .A2(KEYINPUT118), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n537_), .A2(new_n496_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT119), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT119), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n757_), .A2(new_n762_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n497_), .A2(new_n737_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n559_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT57), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n754_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(KEYINPUT57), .A3(new_n559_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n579_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n580_), .A2(new_n677_), .A3(new_n538_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT54), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n439_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n440_), .A2(new_n441_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n537_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(G113gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n732_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n537_), .A2(G113gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n774_), .A2(KEYINPUT59), .A3(new_n775_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n612_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n772_), .B(KEYINPUT54), .Z(new_n782_));
  OAI211_X1 g581(.A(new_n436_), .B(new_n775_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT59), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n779_), .B1(new_n780_), .B2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n732_), .B(new_n777_), .C1(new_n783_), .C2(new_n538_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n778_), .A2(new_n786_), .A3(new_n788_), .ZN(G1340gat));
  AOI21_X1  g588(.A(new_n677_), .B1(new_n780_), .B2(new_n785_), .ZN(new_n790_));
  XOR2_X1   g589(.A(KEYINPUT122), .B(G120gat), .Z(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n677_), .B2(KEYINPUT60), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(KEYINPUT60), .B2(new_n791_), .ZN(new_n793_));
  OAI22_X1  g592(.A1(new_n790_), .A2(new_n791_), .B1(new_n783_), .B2(new_n793_), .ZN(G1341gat));
  AOI21_X1  g593(.A(new_n579_), .B1(new_n780_), .B2(new_n785_), .ZN(new_n795_));
  INV_X1    g594(.A(G127gat), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n612_), .A2(new_n796_), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n795_), .A2(new_n796_), .B1(new_n783_), .B2(new_n797_), .ZN(G1342gat));
  NAND3_X1  g597(.A1(new_n774_), .A2(new_n775_), .A3(new_n585_), .ZN(new_n799_));
  INV_X1    g598(.A(G134gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT123), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n565_), .A2(G134gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n780_), .B2(new_n785_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT123), .B(new_n800_), .C1(new_n783_), .C2(new_n559_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n801_), .A2(new_n803_), .A3(new_n805_), .ZN(G1343gat));
  NOR2_X1   g605(.A1(new_n434_), .A2(new_n253_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n436_), .B(new_n807_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(new_n538_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(new_n266_), .ZN(G1344gat));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n677_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(new_n267_), .ZN(G1345gat));
  NOR2_X1   g611(.A1(new_n808_), .A2(new_n579_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT61), .B(G155gat), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n813_), .B(new_n814_), .Z(G1346gat));
  NOR2_X1   g614(.A1(new_n559_), .A2(G162gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n774_), .A2(new_n807_), .A3(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(G162gat), .B1(new_n808_), .B2(new_n564_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n817_), .A2(new_n818_), .A3(KEYINPUT124), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1347gat));
  NOR2_X1   g622(.A1(new_n441_), .A2(new_n436_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n440_), .B(new_n824_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n825_));
  OAI21_X1  g624(.A(G169gat), .B1(new_n825_), .B2(new_n538_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT125), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT125), .B(G169gat), .C1(new_n825_), .C2(new_n538_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(KEYINPUT62), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n826_), .A2(new_n827_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n825_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n833_), .A2(new_n537_), .A3(new_n390_), .A4(new_n388_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(new_n832_), .A3(new_n834_), .ZN(G1348gat));
  NOR2_X1   g634(.A1(new_n825_), .A2(new_n677_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT126), .B(G176gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n389_), .A2(KEYINPUT126), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n836_), .B2(new_n839_), .ZN(G1349gat));
  NOR2_X1   g639(.A1(new_n825_), .A2(new_n579_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(G183gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n386_), .B2(new_n841_), .ZN(G1350gat));
  OAI21_X1  g642(.A(G190gat), .B1(new_n825_), .B2(new_n564_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n559_), .A2(new_n384_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n825_), .B2(new_n845_), .ZN(G1351gat));
  NAND2_X1  g645(.A1(new_n771_), .A2(new_n773_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n606_), .A2(new_n253_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n824_), .A3(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n538_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n314_), .ZN(G1352gat));
  NOR2_X1   g650(.A1(new_n316_), .A2(KEYINPUT127), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n316_), .A2(KEYINPUT127), .ZN(new_n853_));
  OAI22_X1  g652(.A1(new_n849_), .A2(new_n677_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n849_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n505_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n856_), .B2(new_n852_), .ZN(G1353gat));
  XOR2_X1   g656(.A(KEYINPUT63), .B(G211gat), .Z(new_n858_));
  NAND3_X1  g657(.A1(new_n855_), .A2(new_n612_), .A3(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n849_), .B2(new_n579_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1354gat));
  OAI21_X1  g661(.A(G218gat), .B1(new_n849_), .B2(new_n564_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n559_), .A2(G218gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n849_), .B2(new_n864_), .ZN(G1355gat));
endmodule


