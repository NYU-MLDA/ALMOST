//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT81), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT81), .ZN(new_n205_));
  NOR3_X1   g004(.A1(new_n205_), .A2(G169gat), .A3(G176gat), .ZN(new_n206_));
  OAI211_X1 g005(.A(KEYINPUT24), .B(new_n202_), .C1(new_n204_), .C2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT80), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT26), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT26), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(KEYINPUT80), .A3(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(G183gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n213_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT78), .B1(new_n213_), .B2(KEYINPUT25), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n210_), .B(new_n212_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n213_), .A2(KEYINPUT25), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT79), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n213_), .B2(KEYINPUT25), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n207_), .B1(new_n216_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT82), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n204_), .A2(new_n206_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT82), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n207_), .B(new_n230_), .C1(new_n216_), .C2(new_n221_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n223_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT84), .B(G176gat), .Z(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT83), .B1(new_n234_), .B2(KEYINPUT22), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G169gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n233_), .B(new_n235_), .C1(KEYINPUT83), .C2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n237_), .B(new_n202_), .C1(new_n238_), .C2(new_n226_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G197gat), .B(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G211gat), .A2(G218gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT91), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G211gat), .A2(G218gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n247_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT91), .B1(new_n249_), .B2(new_n244_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT90), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n243_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n241_), .A2(new_n242_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n251_), .B(new_n254_), .C1(new_n252_), .C2(new_n243_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n240_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n202_), .B1(new_n226_), .B2(new_n238_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n236_), .B(KEYINPUT95), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(new_n233_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT25), .B(G183gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT26), .B(G190gat), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n264_), .A2(new_n265_), .B1(new_n228_), .B2(new_n203_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n207_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(new_n226_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n256_), .A2(new_n257_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n260_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G226gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n259_), .A2(new_n271_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT96), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n232_), .A2(new_n270_), .A3(new_n239_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n257_), .B(new_n256_), .C1(new_n263_), .C2(new_n268_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(KEYINPUT20), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n274_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT96), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n259_), .A2(new_n271_), .A3(new_n282_), .A4(new_n275_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G64gat), .B(G92gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT98), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT99), .B(G36gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n289_));
  INV_X1    g088(.A(G8gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n288_), .B(new_n291_), .Z(new_n292_));
  AND2_X1   g091(.A1(new_n292_), .A2(KEYINPUT32), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n284_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n271_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n270_), .B1(new_n232_), .B2(new_n239_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n274_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n278_), .A2(KEYINPUT20), .A3(new_n275_), .A4(new_n279_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n293_), .ZN(new_n300_));
  INV_X1    g099(.A(G155gat), .ZN(new_n301_));
  INV_X1    g100(.A(G162gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G141gat), .ZN(new_n307_));
  INV_X1    g106(.A(G148gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT87), .B1(new_n310_), .B2(new_n316_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(new_n306_), .A4(new_n309_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n313_), .A2(new_n322_), .A3(new_n314_), .ZN(new_n323_));
  OR3_X1    g122(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n309_), .A2(KEYINPUT3), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n303_), .A2(new_n305_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G113gat), .B(G120gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT101), .B1(new_n330_), .B2(new_n334_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n317_), .A2(new_n320_), .B1(new_n328_), .B2(new_n327_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT101), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n333_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT100), .B1(new_n330_), .B2(new_n334_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT100), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n336_), .A2(new_n340_), .A3(new_n333_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n335_), .B(new_n338_), .C1(new_n339_), .C2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  INV_X1    g145(.A(G85gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT0), .B(G57gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT4), .B1(new_n330_), .B2(new_n334_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n342_), .B2(KEYINPUT4), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n345_), .B(new_n351_), .C1(new_n353_), .C2(new_n344_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n344_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n357_));
  AND4_X1   g156(.A1(new_n337_), .A2(new_n321_), .A3(new_n329_), .A4(new_n333_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n337_), .B1(new_n336_), .B2(new_n333_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n330_), .A2(KEYINPUT100), .A3(new_n334_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n340_), .B1(new_n336_), .B2(new_n333_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n357_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n356_), .B1(new_n364_), .B2(new_n352_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n351_), .B1(new_n365_), .B2(new_n345_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n294_), .B(new_n300_), .C1(new_n355_), .C2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT103), .B1(new_n353_), .B2(new_n356_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n343_), .A2(new_n356_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT103), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n370_), .B(new_n344_), .C1(new_n364_), .C2(new_n352_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n368_), .A2(new_n350_), .A3(new_n369_), .A4(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT33), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n354_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n277_), .A2(new_n292_), .A3(new_n281_), .A4(new_n283_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n292_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n284_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .A4(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n342_), .A2(new_n356_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n339_), .A2(new_n341_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n335_), .A2(new_n338_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT4), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n352_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n379_), .B1(new_n384_), .B2(new_n356_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n385_), .A2(KEYINPUT102), .A3(KEYINPUT33), .A4(new_n351_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n365_), .A2(KEYINPUT33), .A3(new_n351_), .A4(new_n345_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT102), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n367_), .B1(new_n378_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G15gat), .B(G43gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT30), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n232_), .A2(new_n396_), .A3(new_n239_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n232_), .B2(new_n239_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n334_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n240_), .A2(KEYINPUT30), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n333_), .A3(new_n397_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G71gat), .B(G99gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n400_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n395_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n400_), .A2(new_n402_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n405_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n400_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n394_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT28), .B(G22gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418_));
  INV_X1    g217(.A(G50gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n336_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n336_), .B2(new_n418_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n417_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n422_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n416_), .A3(new_n420_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n330_), .A2(KEYINPUT29), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT89), .B(G233gat), .Z(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(G228gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n427_), .B(new_n258_), .C1(new_n428_), .C2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n256_), .A2(new_n428_), .A3(new_n257_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n336_), .A2(new_n418_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n433_), .B(new_n430_), .C1(new_n434_), .C2(new_n270_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G78gat), .B(G106gat), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n426_), .B1(new_n438_), .B2(KEYINPUT93), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT93), .ZN(new_n440_));
  INV_X1    g239(.A(new_n437_), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n432_), .A2(new_n435_), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(new_n432_), .B2(new_n435_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n440_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n426_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT92), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n448_), .B(new_n426_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n415_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n391_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n298_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n275_), .B1(new_n259_), .B2(new_n271_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n376_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT104), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT104), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n299_), .A2(new_n457_), .A3(new_n376_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n458_), .A3(new_n375_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT27), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT27), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n377_), .A2(new_n461_), .A3(new_n375_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n355_), .A2(new_n366_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n450_), .A2(new_n414_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n450_), .A2(new_n414_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n463_), .B(new_n464_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n452_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G43gat), .B(G50gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n471_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n469_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT15), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478_));
  INV_X1    g277(.A(G1gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n479_), .B2(new_n290_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G8gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n484_), .B(KEYINPUT75), .Z(new_n485_));
  OR2_X1    g284(.A1(new_n483_), .A2(new_n475_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT76), .Z(new_n488_));
  NAND3_X1  g287(.A1(new_n485_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(KEYINPUT74), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n483_), .A2(new_n475_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(G229gat), .A3(G233gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G169gat), .B(G197gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(new_n307_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT77), .B(G113gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n489_), .A2(new_n493_), .A3(new_n498_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n503_));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT68), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT67), .B(G71gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G78gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT11), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(G78gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n507_), .B(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n506_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n506_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT6), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  OR3_X1    g319(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G85gat), .B(G92gat), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT10), .B(G99gat), .Z(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT66), .B(G106gat), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(KEYINPUT9), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT9), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(G85gat), .A3(G92gat), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n529_), .A2(new_n530_), .A3(new_n532_), .A4(new_n519_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n522_), .A2(KEYINPUT8), .A3(new_n523_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n526_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n517_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n526_), .A2(new_n534_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n533_), .A2(new_n537_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n505_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G230gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n517_), .A2(new_n535_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n539_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT69), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n539_), .A2(KEYINPUT69), .A3(new_n542_), .A4(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n542_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G120gat), .B(G148gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(G204gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT5), .B(G176gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n550_), .A2(new_n552_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n503_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT70), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n558_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n468_), .A2(new_n502_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n477_), .A2(new_n535_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT34), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT35), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n568_), .B(new_n573_), .C1(new_n475_), .C2(new_n535_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n571_), .A2(new_n572_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n575_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n578_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT71), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT71), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n578_), .A2(new_n588_), .A3(new_n584_), .A4(new_n585_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n576_), .A2(new_n583_), .A3(new_n577_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT72), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n483_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n517_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT73), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT16), .B(G183gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT17), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n598_), .B(new_n604_), .Z(new_n605_));
  NOR3_X1   g404(.A1(new_n596_), .A2(KEYINPUT17), .A3(new_n603_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n592_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n567_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n610_), .B2(new_n464_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n586_), .A2(KEYINPUT37), .A3(new_n590_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n591_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(new_n607_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n567_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n464_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n479_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT105), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n621_), .A2(KEYINPUT38), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(KEYINPUT38), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n611_), .B1(new_n622_), .B2(new_n623_), .ZN(G1324gat));
  XNOR2_X1  g423(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n625_));
  INV_X1    g424(.A(new_n463_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n609_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(G8gat), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n628_), .A2(KEYINPUT39), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(KEYINPUT39), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n618_), .A2(new_n290_), .A3(new_n626_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n625_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n632_), .B(new_n625_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n609_), .B2(new_n415_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT41), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n618_), .A2(new_n637_), .A3(new_n415_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n609_), .B2(new_n450_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT42), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n618_), .A2(new_n642_), .A3(new_n450_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1327gat));
  NAND2_X1  g445(.A1(new_n592_), .A2(new_n607_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT109), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n567_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n619_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n468_), .A2(new_n651_), .A3(new_n616_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n468_), .A2(new_n616_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT43), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n468_), .A2(KEYINPUT107), .A3(new_n651_), .A4(new_n616_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n654_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n561_), .A2(new_n565_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n502_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n607_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n659_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n658_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n658_), .B2(new_n662_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n619_), .A2(G29gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n650_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n649_), .A2(new_n670_), .A3(new_n626_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT45), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n658_), .A2(new_n662_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n663_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n658_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n626_), .A3(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(KEYINPUT110), .A3(G36gat), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT110), .B1(new_n676_), .B2(G36gat), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT46), .B(new_n672_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n672_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n679_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n677_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT111), .B(KEYINPUT46), .Z(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1329gat));
  NAND2_X1  g484(.A1(new_n649_), .A2(new_n415_), .ZN(new_n686_));
  INV_X1    g485(.A(G43gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT112), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n665_), .A2(new_n666_), .A3(new_n687_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(new_n415_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n674_), .A2(G43gat), .A3(new_n675_), .A4(new_n415_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(KEYINPUT112), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n688_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT47), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n696_), .B(new_n688_), .C1(new_n691_), .C2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1330gat));
  INV_X1    g497(.A(new_n450_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n665_), .A2(new_n666_), .A3(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT113), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT113), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(G50gat), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n450_), .A2(new_n419_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT114), .Z(new_n705_));
  NAND2_X1  g504(.A1(new_n649_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1331gat));
  NOR2_X1   g506(.A1(new_n566_), .A2(new_n502_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n468_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(new_n617_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n619_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n709_), .A2(new_n608_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n619_), .A2(G57gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n712_), .B2(new_n626_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n710_), .A2(new_n715_), .A3(new_n626_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n712_), .B2(new_n415_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT49), .Z(new_n722_));
  NOR2_X1   g521(.A1(new_n414_), .A2(G71gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT115), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n710_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1334gat));
  AOI21_X1  g525(.A(new_n511_), .B1(new_n712_), .B2(new_n450_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT50), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n710_), .A2(new_n511_), .A3(new_n450_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1335gat));
  AND2_X1   g529(.A1(new_n709_), .A2(new_n648_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n619_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n658_), .A2(new_n607_), .A3(new_n708_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n464_), .A2(new_n347_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(G1336gat));
  AOI21_X1  g534(.A(G92gat), .B1(new_n731_), .B2(new_n626_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n626_), .A2(G92gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT116), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n733_), .B2(new_n738_), .ZN(G1337gat));
  NAND2_X1  g538(.A1(new_n733_), .A2(new_n415_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G99gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n731_), .A2(new_n527_), .A3(new_n415_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g543(.A1(new_n731_), .A2(new_n528_), .A3(new_n450_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n733_), .A2(new_n450_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G106gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT53), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n745_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1339gat));
  INV_X1    g553(.A(new_n466_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT57), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT55), .B1(new_n548_), .B2(new_n549_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n539_), .A2(new_n545_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n551_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n546_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n556_), .B1(new_n757_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT56), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n556_), .C1(new_n757_), .C2(new_n761_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n763_), .A2(new_n502_), .A3(new_n558_), .A4(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n492_), .A2(new_n488_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n485_), .A2(new_n486_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n767_), .B(new_n499_), .C1(new_n768_), .C2(new_n488_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(new_n501_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n770_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n766_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT118), .B(new_n756_), .C1(new_n772_), .C2(new_n592_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n763_), .A2(new_n558_), .A3(new_n770_), .A4(new_n765_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT119), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT58), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(KEYINPUT119), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n616_), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n592_), .B1(new_n766_), .B2(new_n771_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT57), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n773_), .A2(new_n779_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n607_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n615_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n566_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT117), .B1(new_n659_), .B2(new_n785_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(KEYINPUT54), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT117), .B(new_n791_), .C1(new_n659_), .C2(new_n785_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n755_), .B1(new_n784_), .B2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n626_), .A2(new_n464_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(G113gat), .B1(new_n797_), .B2(new_n502_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n795_), .A2(KEYINPUT59), .A3(new_n796_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT59), .B1(new_n795_), .B2(new_n796_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n502_), .A2(G113gat), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT120), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n798_), .B1(new_n803_), .B2(new_n805_), .ZN(G1340gat));
  INV_X1    g605(.A(G120gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n566_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n797_), .B(new_n808_), .C1(KEYINPUT60), .C2(new_n807_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n566_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n807_), .ZN(G1341gat));
  OAI211_X1 g610(.A(G127gat), .B(new_n661_), .C1(new_n799_), .C2(new_n801_), .ZN(new_n812_));
  INV_X1    g611(.A(G127gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n795_), .A2(new_n796_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n607_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT121), .B(new_n813_), .C1(new_n814_), .C2(new_n607_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n812_), .A2(new_n817_), .A3(new_n818_), .ZN(G1342gat));
  AOI21_X1  g618(.A(G134gat), .B1(new_n797_), .B2(new_n592_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n615_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g621(.A1(new_n784_), .A2(new_n794_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n796_), .A2(new_n465_), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(KEYINPUT122), .Z(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n660_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(new_n307_), .ZN(G1344gat));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n566_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(new_n308_), .ZN(G1345gat));
  INV_X1    g629(.A(new_n826_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n301_), .A3(new_n661_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G155gat), .B1(new_n826_), .B2(new_n607_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n832_), .A2(new_n835_), .A3(new_n833_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(G1346gat));
  NOR3_X1   g638(.A1(new_n826_), .A2(new_n302_), .A3(new_n615_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n831_), .A2(new_n592_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n302_), .B2(new_n841_), .ZN(G1347gat));
  NOR2_X1   g641(.A1(new_n463_), .A2(new_n619_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n415_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n823_), .A2(new_n502_), .A3(new_n699_), .A4(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n450_), .B1(new_n784_), .B2(new_n794_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n849_), .A2(KEYINPUT124), .A3(new_n502_), .A4(new_n845_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n850_), .A3(G169gat), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n823_), .A2(new_n699_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n844_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n502_), .A3(new_n262_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n848_), .A2(new_n850_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n853_), .A2(new_n856_), .A3(new_n857_), .ZN(G1348gat));
  OR2_X1    g657(.A1(new_n854_), .A2(KEYINPUT125), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n854_), .A2(KEYINPUT125), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n659_), .A2(G176gat), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n859_), .A2(new_n845_), .A3(new_n860_), .A4(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n855_), .A2(new_n659_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n233_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1349gat));
  NAND4_X1  g664(.A1(new_n859_), .A2(new_n661_), .A3(new_n845_), .A4(new_n860_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n607_), .A2(new_n264_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n866_), .A2(new_n213_), .B1(new_n855_), .B2(new_n867_), .ZN(G1350gat));
  NAND3_X1  g667(.A1(new_n855_), .A2(new_n265_), .A3(new_n592_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n854_), .A2(new_n615_), .A3(new_n844_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n209_), .ZN(G1351gat));
  AND3_X1   g670(.A1(new_n823_), .A2(new_n465_), .A3(new_n843_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n502_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g673(.A(G204gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT126), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT126), .B(G204gat), .Z(new_n877_));
  NAND3_X1  g676(.A1(new_n823_), .A2(new_n465_), .A3(new_n843_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n566_), .ZN(new_n879_));
  MUX2_X1   g678(.A(new_n876_), .B(new_n877_), .S(new_n879_), .Z(G1353gat));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  AND2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  NOR4_X1   g681(.A1(new_n878_), .A2(new_n607_), .A3(new_n881_), .A4(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n872_), .A2(new_n661_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n881_), .ZN(G1354gat));
  NAND3_X1  g684(.A1(new_n872_), .A2(KEYINPUT127), .A3(new_n592_), .ZN(new_n886_));
  INV_X1    g685(.A(G218gat), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n878_), .B2(new_n591_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n887_), .A3(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n872_), .A2(G218gat), .A3(new_n616_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1355gat));
endmodule


