//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT85), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n202_), .A2(new_n203_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT30), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT23), .ZN(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G190gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT81), .B(G190gat), .Z(new_n221_));
  OAI211_X1 g020(.A(new_n218_), .B(new_n220_), .C1(new_n221_), .C2(new_n219_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n215_), .A2(KEYINPUT24), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT82), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(KEYINPUT82), .A3(new_n224_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n217_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n221_), .A2(G183gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n230_), .A2(new_n212_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(new_n213_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n210_), .B1(new_n229_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n234_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n217_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n228_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT82), .B1(new_n222_), .B2(new_n224_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n240_), .A3(KEYINPUT30), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT84), .B(G15gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n235_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n209_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n235_), .A2(new_n241_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n244_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n235_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n208_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G71gat), .B(G99gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT83), .B(G43gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT31), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n248_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n248_), .B2(new_n252_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT86), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT86), .A3(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n264_), .A2(new_n266_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT1), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(G155gat), .A3(G162gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n261_), .A2(new_n267_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n271_), .A2(new_n275_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT28), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(new_n285_), .A3(new_n282_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G22gat), .B(G50gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT89), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n286_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n287_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT89), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n288_), .ZN(new_n296_));
  INV_X1    g095(.A(G197gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT87), .B1(new_n297_), .B2(G204gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299_));
  INV_X1    g098(.A(G204gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(G197gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT21), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(G204gat), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n298_), .A2(new_n301_), .A3(new_n302_), .A4(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n297_), .A2(G204gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n300_), .A2(G197gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT21), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n298_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n308_), .A2(new_n302_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n311_), .A2(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n281_), .A2(new_n282_), .ZN(new_n316_));
  OAI211_X1 g115(.A(G228gat), .B(G233gat), .C1(new_n315_), .C2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n312_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n313_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G228gat), .A2(G233gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n316_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n291_), .A2(new_n296_), .A3(new_n317_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n323_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n294_), .A2(new_n288_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(KEYINPUT89), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G78gat), .B(G106gat), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n324_), .A2(new_n329_), .A3(new_n327_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n260_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n336_), .A2(KEYINPUT33), .ZN(new_n337_));
  INV_X1    g136(.A(new_n281_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n208_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n202_), .A2(new_n203_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n281_), .B1(new_n207_), .B2(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(KEYINPUT4), .A3(new_n341_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT94), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n339_), .A2(new_n348_), .A3(KEYINPUT4), .A4(new_n341_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n339_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n349_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n345_), .B1(new_n353_), .B2(new_n344_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT0), .B(G57gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n337_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n337_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n346_), .A2(KEYINPUT94), .B1(new_n350_), .B2(new_n351_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n343_), .B1(new_n362_), .B2(new_n349_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n358_), .B(new_n361_), .C1(new_n363_), .C2(new_n345_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n343_), .B1(new_n342_), .B2(KEYINPUT96), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(KEYINPUT96), .B2(new_n342_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n366_), .B(new_n359_), .C1(new_n344_), .C2(new_n353_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n360_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT18), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n370_), .B(new_n371_), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT19), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n229_), .A2(new_n234_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(new_n315_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT26), .B(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n218_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n237_), .A2(KEYINPUT90), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT90), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n217_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n224_), .B(new_n381_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G169gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT91), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n214_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n212_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n388_), .B(new_n223_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n320_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n376_), .B1(new_n379_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n320_), .B1(new_n229_), .B2(new_n234_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n315_), .A2(new_n385_), .A3(new_n391_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n395_), .A2(KEYINPUT20), .A3(new_n396_), .A4(new_n376_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n373_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT92), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n236_), .A2(new_n240_), .A3(new_n315_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n393_), .A2(KEYINPUT20), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n375_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n372_), .A3(new_n397_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n399_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT93), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT92), .B(new_n373_), .C1(new_n394_), .C2(new_n398_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n406_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n368_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n402_), .A2(new_n375_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n395_), .A2(KEYINPUT20), .A3(new_n396_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n375_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT97), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n372_), .A2(KEYINPUT32), .ZN(new_n415_));
  OR3_X1    g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n354_), .A2(new_n359_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n358_), .B1(new_n363_), .B2(new_n345_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n403_), .A2(new_n397_), .A3(new_n415_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n414_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n335_), .B1(new_n410_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n332_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n329_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n425_));
  OAI22_X1  g224(.A1(new_n257_), .A2(new_n258_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n256_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n246_), .A2(new_n247_), .A3(new_n209_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n208_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n248_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n430_), .A2(new_n331_), .A3(new_n332_), .A4(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n419_), .B1(new_n426_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT27), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n405_), .A2(new_n434_), .A3(new_n407_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT27), .B(new_n404_), .C1(new_n413_), .C2(new_n372_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n423_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT73), .B(G1gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G190gat), .B(G218gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT71), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G134gat), .B(G162gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT69), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT65), .ZN(new_n448_));
  OAI22_X1  g247(.A1(new_n448_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT7), .ZN(new_n450_));
  INV_X1    g249(.A(G99gat), .ZN(new_n451_));
  INV_X1    g250(.A(G106gat), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .A4(KEYINPUT65), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(G99gat), .B2(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n449_), .B(new_n453_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G85gat), .ZN(new_n459_));
  INV_X1    g258(.A(G92gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT8), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT8), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n458_), .A2(new_n466_), .A3(new_n463_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT64), .ZN(new_n468_));
  INV_X1    g267(.A(new_n462_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(KEYINPUT9), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT9), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n462_), .A2(KEYINPUT64), .A3(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n470_), .A2(new_n472_), .A3(new_n473_), .A4(new_n461_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n455_), .A2(new_n457_), .ZN(new_n475_));
  OR2_X1    g274(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n476_), .A2(new_n452_), .A3(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n465_), .A2(new_n467_), .B1(new_n474_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G29gat), .B(G36gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G43gat), .B(G50gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n482_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT15), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(KEYINPUT15), .A3(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n447_), .B1(new_n480_), .B2(new_n489_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n483_), .A2(KEYINPUT15), .A3(new_n484_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT15), .B1(new_n483_), .B2(new_n484_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n479_), .A2(new_n474_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n458_), .A2(new_n466_), .A3(new_n463_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n466_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n497_), .A3(KEYINPUT69), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n480_), .A2(new_n485_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n490_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT68), .B(KEYINPUT35), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n446_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n490_), .A2(KEYINPUT70), .A3(new_n498_), .A4(new_n499_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G232gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n501_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n493_), .A2(new_n497_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n509_), .A2(new_n447_), .B1(new_n485_), .B2(new_n480_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n507_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n510_), .A2(KEYINPUT70), .A3(new_n498_), .A4(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n502_), .A2(new_n508_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n444_), .A2(new_n445_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n502_), .A2(new_n508_), .A3(new_n512_), .A4(new_n514_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n517_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT72), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT79), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G57gat), .B(G64gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G71gat), .B(G78gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(KEYINPUT11), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(KEYINPUT11), .ZN(new_n529_));
  INV_X1    g328(.A(new_n527_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n526_), .A2(KEYINPUT11), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n528_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G231gat), .ZN(new_n534_));
  INV_X1    g333(.A(G233gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n528_), .B(new_n537_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G1gat), .B(G8gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT74), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543_));
  INV_X1    g342(.A(G8gat), .ZN(new_n544_));
  INV_X1    g343(.A(G1gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT73), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(G1gat), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n544_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n542_), .B(new_n543_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(new_n440_), .B2(new_n544_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n542_), .B1(new_n553_), .B2(new_n543_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n541_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n549_), .A2(new_n550_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n543_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT74), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(new_n551_), .A3(new_n540_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n539_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n536_), .A2(new_n555_), .A3(new_n559_), .A4(new_n538_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT75), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT75), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(new_n565_), .A3(new_n562_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n568_));
  XOR2_X1   g367(.A(G183gat), .B(G211gat), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G127gat), .B(G155gat), .Z(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n569_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n568_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n574_), .A3(new_n568_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n567_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n564_), .A2(new_n566_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT17), .B1(new_n580_), .B2(new_n575_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n576_), .A2(new_n567_), .A3(new_n577_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT77), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n581_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT77), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n563_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT78), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n579_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n579_), .B2(new_n587_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n525_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n579_), .A2(new_n587_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT78), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n579_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(KEYINPUT79), .A3(new_n594_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n520_), .A2(new_n524_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT80), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n555_), .A2(new_n559_), .A3(new_n485_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n485_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n560_), .A2(new_n493_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n555_), .A2(new_n559_), .A3(new_n485_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n598_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G113gat), .B(G141gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G169gat), .B(G197gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n607_), .B(new_n608_), .Z(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n597_), .B1(new_n606_), .B2(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n602_), .A2(new_n605_), .A3(KEYINPUT80), .A4(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n606_), .A2(new_n610_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n533_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n497_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n533_), .B(new_n494_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n617_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(KEYINPUT12), .A3(new_n620_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT12), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n497_), .A2(new_n623_), .A3(new_n618_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n621_), .B1(new_n625_), .B2(new_n617_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT5), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n630_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n617_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n632_), .B1(new_n634_), .B2(new_n621_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n631_), .A2(KEYINPUT66), .A3(new_n635_), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n626_), .A2(KEYINPUT66), .A3(new_n630_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT13), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n637_), .A3(KEYINPUT13), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n596_), .A2(new_n616_), .A3(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n439_), .A2(new_n419_), .A3(new_n440_), .A4(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT38), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n423_), .A2(new_n438_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n521_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n642_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n615_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n593_), .A2(new_n594_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n646_), .A2(new_n647_), .A3(new_n652_), .ZN(new_n653_));
  AOI211_X1 g452(.A(KEYINPUT98), .B(new_n545_), .C1(new_n653_), .C2(new_n419_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n419_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(G1gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n645_), .B1(new_n654_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT99), .ZN(G1324gat));
  AND2_X1   g458(.A1(new_n439_), .A2(new_n643_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n435_), .A2(new_n436_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n544_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n653_), .A2(new_n661_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(G8gat), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT39), .B(new_n544_), .C1(new_n653_), .C2(new_n661_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g467(.A1(new_n653_), .A2(new_n259_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n669_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(new_n669_), .B2(G15gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n660_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n260_), .A2(G15gat), .ZN(new_n673_));
  OAI22_X1  g472(.A1(new_n670_), .A2(new_n671_), .B1(new_n672_), .B2(new_n673_), .ZN(G1326gat));
  OR3_X1    g473(.A1(new_n672_), .A2(G22gat), .A3(new_n334_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n653_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G22gat), .B1(new_n676_), .B2(new_n334_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n677_), .A2(KEYINPUT101), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(KEYINPUT101), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n675_), .B1(new_n681_), .B2(new_n682_), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n524_), .A2(new_n520_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(new_n423_), .B2(new_n438_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n591_), .A2(new_n595_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT43), .B(new_n685_), .C1(new_n423_), .C2(new_n438_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n688_), .A2(new_n649_), .A3(new_n690_), .A4(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n689_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n695_), .A2(KEYINPUT44), .A3(new_n649_), .A4(new_n691_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n694_), .A2(G29gat), .A3(new_n419_), .A4(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(G29gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n689_), .A2(new_n521_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n439_), .A2(KEYINPUT102), .A3(new_n649_), .A4(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n699_), .B(new_n649_), .C1(new_n423_), .C2(new_n438_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n419_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n697_), .A2(new_n706_), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n694_), .A2(new_n661_), .A3(new_n696_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G36gat), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n437_), .A2(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n700_), .A2(new_n703_), .A3(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT45), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(new_n712_), .A3(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n694_), .A2(G43gat), .A3(new_n259_), .A4(new_n696_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n700_), .A2(new_n259_), .A3(new_n703_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT103), .B(G43gat), .Z(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(KEYINPUT104), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT104), .B1(new_n719_), .B2(new_n720_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT47), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n718_), .B(new_n725_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  NAND4_X1  g526(.A1(new_n694_), .A2(G50gat), .A3(new_n333_), .A4(new_n696_), .ZN(new_n728_));
  INV_X1    g527(.A(G50gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n729_), .B1(new_n704_), .B2(new_n334_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n648_), .A2(new_n596_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT105), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n439_), .A3(new_n615_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n735_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n705_), .A2(G57gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n646_), .A2(new_n647_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n690_), .A2(new_n642_), .A3(new_n616_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n705_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n739_), .A2(new_n743_), .ZN(G1332gat));
  NOR2_X1   g543(.A1(new_n437_), .A2(G64gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n736_), .A2(new_n737_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G64gat), .B1(new_n742_), .B2(new_n437_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(KEYINPUT48), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(KEYINPUT48), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n748_), .B2(new_n749_), .ZN(G1333gat));
  NOR2_X1   g549(.A1(new_n260_), .A2(G71gat), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT107), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n736_), .A2(new_n737_), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G71gat), .B1(new_n742_), .B2(new_n260_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(KEYINPUT49), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(KEYINPUT49), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(G1334gat));
  NOR2_X1   g556(.A1(new_n334_), .A2(G78gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n736_), .A2(new_n737_), .A3(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G78gat), .B1(new_n742_), .B2(new_n334_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(KEYINPUT50), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(KEYINPUT50), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n642_), .A2(new_n616_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n695_), .A2(new_n691_), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n705_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n439_), .A2(new_n699_), .A3(new_n764_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n459_), .A3(new_n419_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1336gat));
  OAI21_X1  g568(.A(G92gat), .B1(new_n765_), .B2(new_n437_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n460_), .A3(new_n661_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT108), .Z(G1337gat));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(KEYINPUT51), .ZN(new_n775_));
  OAI21_X1  g574(.A(G99gat), .B1(new_n765_), .B2(new_n260_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n767_), .A2(new_n476_), .A3(new_n477_), .A4(new_n259_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n774_), .A2(KEYINPUT51), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1338gat));
  OAI21_X1  g579(.A(G106gat), .B1(new_n765_), .B2(new_n334_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  XOR2_X1   g582(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n784_));
  OAI211_X1 g583(.A(G106gat), .B(new_n784_), .C1(new_n765_), .C2(new_n334_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n767_), .A2(new_n452_), .A3(new_n333_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n783_), .A2(new_n789_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1339gat));
  NAND4_X1  g590(.A1(new_n642_), .A2(new_n684_), .A3(new_n615_), .A4(new_n689_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT54), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n596_), .A2(new_n794_), .A3(new_n615_), .A4(new_n642_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n622_), .A2(new_n633_), .A3(new_n624_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n799_), .A2(new_n634_), .A3(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n625_), .A2(new_n800_), .A3(new_n617_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n632_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n798_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n630_), .B1(new_n634_), .B2(new_n800_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n625_), .A2(new_n617_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT55), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT56), .B(new_n806_), .C1(new_n808_), .C2(new_n799_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(new_n805_), .A3(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT113), .B(new_n798_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n598_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n603_), .A2(new_n604_), .A3(new_n599_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n610_), .ZN(new_n814_));
  AOI221_X4 g613(.A(new_n814_), .B1(new_n626_), .B2(new_n630_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n810_), .A2(new_n811_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n684_), .B1(new_n797_), .B2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n810_), .A2(new_n815_), .A3(KEYINPUT58), .A4(new_n811_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n804_), .A2(KEYINPUT111), .A3(new_n809_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n613_), .A2(new_n614_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n801_), .A2(new_n803_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(KEYINPUT56), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(new_n820_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n814_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n647_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n817_), .A2(new_n818_), .B1(new_n827_), .B2(KEYINPUT57), .ZN(new_n828_));
  INV_X1    g627(.A(new_n827_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(KEYINPUT112), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n827_), .B2(KEYINPUT57), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n828_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n796_), .B1(new_n834_), .B2(new_n650_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n661_), .A2(new_n705_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n432_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n616_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT59), .B1(new_n835_), .B2(new_n838_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n824_), .A2(new_n826_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(KEYINPUT57), .A3(new_n521_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n816_), .A2(new_n797_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n685_), .A3(new_n818_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n827_), .A2(KEYINPUT57), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n690_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n793_), .A2(new_n795_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n838_), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n841_), .A2(KEYINPUT114), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT114), .B1(new_n841_), .B2(new_n852_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(G113gat), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n616_), .A2(KEYINPUT115), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(G113gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n840_), .B1(new_n855_), .B2(new_n859_), .ZN(G1340gat));
  NAND3_X1  g659(.A1(new_n841_), .A2(new_n648_), .A3(new_n852_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G120gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n642_), .A2(KEYINPUT60), .ZN(new_n863_));
  MUX2_X1   g662(.A(new_n863_), .B(KEYINPUT60), .S(G120gat), .Z(new_n864_));
  NAND2_X1  g663(.A1(new_n839_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1341gat));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n839_), .A2(new_n867_), .A3(new_n689_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n853_), .A2(new_n854_), .A3(new_n650_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1342gat));
  INV_X1    g669(.A(G134gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n839_), .A2(new_n871_), .A3(new_n647_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n853_), .A2(new_n854_), .A3(new_n684_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n871_), .ZN(G1343gat));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875_));
  INV_X1    g674(.A(new_n426_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n836_), .A2(new_n876_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n877_), .A2(KEYINPUT116), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(KEYINPUT116), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n835_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n875_), .B1(new_n881_), .B2(new_n616_), .ZN(new_n882_));
  NOR4_X1   g681(.A1(new_n835_), .A2(new_n880_), .A3(KEYINPUT118), .A4(new_n615_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT117), .B(G141gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1344gat));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n648_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT119), .B(G148gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1345gat));
  NAND2_X1  g688(.A1(new_n881_), .A2(new_n689_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n881_), .B2(new_n647_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n685_), .A2(G162gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT120), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n881_), .B2(new_n895_), .ZN(G1347gat));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897_));
  INV_X1    g696(.A(new_n847_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n828_), .A2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n796_), .B1(new_n899_), .B2(new_n690_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n661_), .A2(new_n705_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n432_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n897_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n850_), .A2(KEYINPUT122), .A3(new_n902_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n904_), .A2(new_n387_), .A3(new_n616_), .A4(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n902_), .A2(new_n616_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n689_), .B1(new_n828_), .B2(new_n898_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT121), .B(new_n908_), .C1(new_n909_), .C2(new_n796_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G169gat), .ZN(new_n911_));
  AOI21_X1  g710(.A(KEYINPUT121), .B1(new_n850_), .B2(new_n908_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n911_), .A2(new_n912_), .A3(KEYINPUT62), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n907_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n213_), .B1(new_n915_), .B2(KEYINPUT121), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n900_), .B2(new_n907_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n914_), .B1(new_n916_), .B2(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n906_), .B1(new_n913_), .B2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT123), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n922_), .B(new_n906_), .C1(new_n913_), .C2(new_n919_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1348gat));
  NAND2_X1  g723(.A1(new_n904_), .A2(new_n905_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n214_), .B1(new_n925_), .B2(new_n642_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n835_), .A2(new_n333_), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n901_), .A2(new_n214_), .A3(new_n260_), .A4(new_n642_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n926_), .A2(KEYINPUT124), .A3(new_n929_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1349gat));
  NOR2_X1   g733(.A1(new_n650_), .A2(new_n218_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT125), .B1(new_n925_), .B2(new_n936_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n901_), .A2(new_n260_), .A3(new_n690_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n927_), .A2(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n937_), .B1(G183gat), .B2(new_n939_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n925_), .A2(KEYINPUT125), .A3(new_n936_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n925_), .B2(new_n684_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n647_), .A2(new_n380_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n925_), .B2(new_n944_), .ZN(G1351gat));
  NOR3_X1   g744(.A1(new_n835_), .A2(new_n426_), .A3(new_n901_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n616_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n297_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(KEYINPUT126), .B(G197gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n947_), .B2(new_n950_), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n946_), .A2(new_n648_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g752(.A1(new_n946_), .A2(new_n651_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AND2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n954_), .A2(new_n955_), .A3(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n957_), .B1(new_n954_), .B2(new_n955_), .ZN(G1354gat));
  INV_X1    g757(.A(G218gat), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n946_), .A2(new_n959_), .A3(new_n647_), .ZN(new_n960_));
  AND2_X1   g759(.A1(new_n946_), .A2(new_n685_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n961_), .B2(new_n959_), .ZN(G1355gat));
endmodule


