//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT6), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT7), .ZN(new_n205_));
  INV_X1    g004(.A(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n202_), .B1(new_n204_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n203_), .B(KEYINPUT6), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n212_), .A2(KEYINPUT67), .A3(new_n208_), .A4(new_n209_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  XOR2_X1   g013(.A(G85gat), .B(G92gat), .Z(new_n215_));
  NAND4_X1  g014(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n210_), .B1(new_n212_), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(new_n212_), .B2(new_n217_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n219_), .A2(new_n215_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n216_), .B1(new_n220_), .B2(new_n214_), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n204_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n225_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n215_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT10), .B(G99gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT65), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n226_), .B(new_n229_), .C1(new_n231_), .C2(G106gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G78gat), .Z(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n235_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n221_), .A2(new_n232_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT12), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n221_), .B2(new_n232_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G230gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT64), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n248_), .B(new_n216_), .C1(new_n220_), .C2(new_n214_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n214_), .B1(new_n219_), .B2(new_n215_), .ZN(new_n250_));
  AND4_X1   g049(.A1(new_n214_), .A2(new_n211_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT71), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n252_), .A3(new_n232_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n236_), .B(KEYINPUT12), .C1(new_n237_), .C2(new_n238_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT72), .B1(new_n253_), .B2(new_n255_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n244_), .B(new_n247_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n243_), .A2(KEYINPUT70), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n240_), .B1(new_n242_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n246_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G120gat), .B(G148gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(new_n264_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n275_), .A2(KEYINPUT13), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT13), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n271_), .A2(new_n275_), .A3(KEYINPUT13), .A4(new_n273_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT75), .ZN(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT80), .B(G1gat), .Z(new_n282_));
  INV_X1    g081(.A(G8gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT14), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G1gat), .B(G8gat), .Z(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G29gat), .B(G36gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(G43gat), .B(G50gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT84), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n290_), .B(new_n294_), .Z(new_n295_));
  NAND2_X1  g094(.A1(G229gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n290_), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n293_), .B(KEYINPUT15), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n290_), .A2(new_n294_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n296_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G113gat), .B(G141gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G169gat), .B(G197gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n305_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n278_), .A2(new_n311_), .A3(new_n279_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n281_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G231gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n239_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(new_n299_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G127gat), .B(G155gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(G183gat), .B(G211gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(KEYINPUT17), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(KEYINPUT17), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT83), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n316_), .A2(KEYINPUT82), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n313_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G113gat), .B(G120gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G169gat), .ZN(new_n334_));
  INV_X1    g133(.A(G176gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT85), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT85), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT23), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(G183gat), .A3(G190gat), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n336_), .B(new_n341_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT86), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n338_), .A4(new_n340_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n352_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n351_), .B1(new_n341_), .B2(new_n350_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n348_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT87), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n338_), .A2(new_n340_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT86), .B1(new_n363_), .B2(new_n349_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n364_), .A2(new_n352_), .A3(new_n357_), .A4(new_n354_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT87), .A3(new_n348_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT30), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G71gat), .B(G99gat), .ZN(new_n369_));
  INV_X1    g168(.A(G43gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G15gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n371_), .B(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n368_), .A2(new_n374_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT31), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n375_), .A2(new_n376_), .A3(KEYINPUT31), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n333_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n332_), .A3(new_n377_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383_));
  INV_X1    g182(.A(G141gat), .ZN(new_n384_));
  INV_X1    g183(.A(G148gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT2), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n386_), .B(new_n387_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n388_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT90), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n387_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G141gat), .A2(G148gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT2), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n396_), .A2(new_n397_), .A3(new_n391_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n393_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT88), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n384_), .A2(new_n385_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n398_), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n406_), .B(KEYINPUT1), .Z(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n412_), .B2(new_n405_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n409_), .A2(new_n414_), .A3(new_n332_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n407_), .B1(new_n393_), .B2(new_n402_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n333_), .B1(new_n416_), .B2(new_n413_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(new_n333_), .C1(new_n416_), .C2(new_n413_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT97), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n415_), .A2(KEYINPUT4), .A3(new_n417_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n418_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n419_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT0), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G57gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(new_n222_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n431_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n433_), .B(new_n419_), .C1(new_n422_), .C2(new_n425_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n380_), .A2(new_n382_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT19), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n350_), .A2(new_n337_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT95), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n357_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n357_), .B2(new_n441_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n354_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n348_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT91), .B(G197gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(G204gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT21), .ZN(new_n449_));
  INV_X1    g248(.A(G197gat), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n448_), .B(new_n449_), .C1(new_n450_), .C2(G204gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(G211gat), .B(G218gat), .Z(new_n452_));
  INV_X1    g251(.A(G204gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n449_), .B1(G197gat), .B2(G204gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n452_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n451_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n448_), .B1(new_n450_), .B2(G204gat), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n452_), .A2(KEYINPUT21), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT20), .B1(new_n446_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT96), .B1(new_n367_), .B2(new_n461_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT96), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n451_), .A2(new_n456_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n466_));
  AOI211_X1 g265(.A(new_n465_), .B(new_n466_), .C1(new_n362_), .C2(new_n366_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n440_), .B(new_n463_), .C1(new_n464_), .C2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n446_), .B2(new_n461_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n362_), .A2(new_n366_), .A3(new_n466_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n440_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G8gat), .B(G36gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT18), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G64gat), .B(G92gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n468_), .A2(new_n473_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT27), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n365_), .A2(KEYINPUT87), .A3(new_n348_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT87), .B1(new_n365_), .B2(new_n348_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n461_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n465_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n367_), .A2(KEYINPUT96), .A3(new_n461_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n462_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n472_), .B1(new_n489_), .B2(new_n440_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n483_), .B1(new_n490_), .B2(new_n480_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n439_), .B(new_n463_), .C1(new_n464_), .C2(new_n467_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n470_), .A2(new_n471_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n440_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n478_), .A3(new_n494_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n482_), .A2(new_n483_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n416_), .B2(new_n413_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n461_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G228gat), .A2(G233gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n416_), .A2(new_n413_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n500_), .B(new_n461_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G78gat), .B(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n502_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT93), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n502_), .A2(KEYINPUT93), .A3(new_n505_), .A4(new_n507_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n461_), .A2(new_n500_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n409_), .A2(new_n414_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(KEYINPUT29), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n500_), .B1(new_n498_), .B2(new_n461_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n506_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n510_), .A2(new_n511_), .A3(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT28), .B1(new_n513_), .B2(KEYINPUT29), .ZN(new_n518_));
  NOR4_X1   g317(.A1(new_n416_), .A2(KEYINPUT28), .A3(KEYINPUT29), .A4(new_n413_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G22gat), .B(G50gat), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n521_), .B1(new_n525_), .B2(new_n519_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n517_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n516_), .A2(new_n508_), .A3(new_n523_), .A4(new_n526_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n527_), .A2(KEYINPUT94), .A3(new_n508_), .A4(new_n516_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n496_), .A2(KEYINPUT101), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT101), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n468_), .A2(new_n473_), .A3(new_n480_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n480_), .B1(new_n468_), .B2(new_n473_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n483_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n481_), .A2(new_n495_), .A3(KEYINPUT27), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n537_), .B1(new_n542_), .B2(new_n534_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n437_), .B1(new_n536_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n492_), .A2(new_n546_), .A3(new_n494_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT98), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT98), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n492_), .A2(new_n549_), .A3(new_n546_), .A4(new_n494_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n468_), .A2(new_n473_), .A3(new_n545_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n435_), .A2(new_n548_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT33), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n421_), .B(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(new_n418_), .A3(new_n423_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n415_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n431_), .A2(new_n557_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n434_), .A2(new_n553_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(new_n424_), .A3(new_n423_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n560_), .A2(KEYINPUT33), .A3(new_n419_), .A4(new_n433_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n559_), .A2(new_n481_), .A3(new_n479_), .A4(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n552_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n535_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT99), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n534_), .B1(new_n562_), .B2(new_n552_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n532_), .A2(new_n533_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n507_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n509_), .B2(new_n508_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n527_), .B1(new_n571_), .B2(new_n511_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n436_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT100), .B1(new_n573_), .B2(new_n542_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n496_), .A2(new_n575_), .A3(new_n436_), .A4(new_n534_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n565_), .A2(new_n568_), .A3(new_n574_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n380_), .A2(new_n382_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n544_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT77), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n221_), .A2(new_n232_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT34), .ZN(new_n583_));
  OAI22_X1  g382(.A1(new_n581_), .A2(new_n293_), .B1(KEYINPUT35), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n583_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT35), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n253_), .A2(new_n300_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n580_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n588_), .A2(new_n580_), .A3(new_n589_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G190gat), .B(G218gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(KEYINPUT36), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n584_), .A2(KEYINPUT76), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n589_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n584_), .A2(KEYINPUT76), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n587_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n593_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n596_), .B(KEYINPUT36), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT78), .Z(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n579_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n329_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G1gat), .B1(new_n612_), .B2(new_n436_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n313_), .A2(new_n579_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n606_), .B(KEYINPUT79), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n604_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n615_), .B1(new_n619_), .B2(new_n603_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n603_), .A2(new_n615_), .A3(new_n607_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(new_n328_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n614_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n435_), .A2(new_n282_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n613_), .B1(new_n630_), .B2(new_n631_), .ZN(G1324gat));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n283_), .A3(new_n542_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n611_), .A2(new_n542_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G8gat), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(KEYINPUT39), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(KEYINPUT39), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g438(.A(G15gat), .B1(new_n612_), .B2(new_n578_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT41), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(KEYINPUT41), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n625_), .A2(G15gat), .A3(new_n578_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n641_), .A2(new_n642_), .A3(new_n643_), .ZN(G1326gat));
  OAI21_X1  g443(.A(G22gat), .B1(new_n612_), .B2(new_n535_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT42), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n535_), .A2(G22gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n625_), .B2(new_n647_), .ZN(G1327gat));
  XOR2_X1   g447(.A(new_n326_), .B(new_n327_), .Z(new_n649_));
  OR3_X1    g448(.A1(new_n649_), .A2(new_n608_), .A3(KEYINPUT104), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT104), .B1(new_n649_), .B2(new_n608_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n614_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G29gat), .B1(new_n654_), .B2(new_n435_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n576_), .B(new_n574_), .C1(new_n567_), .C2(new_n566_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n568_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n578_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n544_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n623_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n603_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT37), .B1(new_n663_), .B2(new_n618_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n621_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n579_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n313_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n667_), .A2(KEYINPUT44), .A3(new_n668_), .A4(new_n328_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n669_), .A2(G29gat), .A3(new_n435_), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n313_), .B(new_n649_), .C1(new_n662_), .C2(new_n666_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n655_), .B1(new_n670_), .B2(new_n674_), .ZN(G1328gat));
  OR2_X1    g474(.A1(new_n496_), .A2(KEYINPUT106), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n496_), .A2(KEYINPUT106), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n653_), .A2(G36gat), .A3(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT45), .Z(new_n681_));
  OAI211_X1 g480(.A(new_n669_), .B(new_n542_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT105), .B1(new_n682_), .B2(G36gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT46), .B(new_n681_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  INV_X1    g488(.A(new_n578_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n674_), .A2(G43gat), .A3(new_n690_), .A4(new_n669_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n370_), .B1(new_n653_), .B2(new_n578_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g493(.A(G50gat), .B1(new_n654_), .B2(new_n534_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n669_), .A2(G50gat), .A3(new_n534_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n674_), .ZN(G1331gat));
  NAND2_X1  g496(.A1(new_n281_), .A2(new_n312_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n328_), .A2(new_n310_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n610_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(G57gat), .A3(new_n435_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n310_), .B1(new_n281_), .B2(new_n312_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n624_), .A2(new_n660_), .A3(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n436_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n706_), .B2(G57gat), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT107), .Z(G1332gat));
  OR3_X1    g507(.A1(new_n705_), .A2(G64gat), .A3(new_n679_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n702_), .A2(new_n678_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(G64gat), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G64gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT109), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n701_), .B2(new_n578_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT49), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n578_), .A2(G71gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n705_), .B2(new_n718_), .ZN(G1334gat));
  OR3_X1    g518(.A1(new_n705_), .A2(G78gat), .A3(new_n535_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G78gat), .B1(new_n701_), .B2(new_n535_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(KEYINPUT50), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(KEYINPUT50), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(G1335gat));
  NAND3_X1  g523(.A1(new_n667_), .A2(new_n328_), .A3(new_n704_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n436_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n652_), .A2(new_n704_), .A3(new_n660_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT110), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n652_), .A2(new_n704_), .A3(new_n729_), .A4(new_n660_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(new_n222_), .A3(new_n435_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n726_), .A2(new_n732_), .ZN(G1336gat));
  OAI21_X1  g532(.A(G92gat), .B1(new_n725_), .B2(new_n679_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n223_), .A3(new_n542_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1337gat));
  NOR2_X1   g535(.A1(new_n578_), .A2(new_n231_), .ZN(new_n737_));
  AOI22_X1  g536(.A1(new_n731_), .A2(new_n737_), .B1(KEYINPUT112), .B2(KEYINPUT51), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n667_), .A2(new_n690_), .A3(new_n328_), .A4(new_n704_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(new_n740_), .A3(G99gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n739_), .B2(G99gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT113), .ZN(new_n744_));
  NOR2_X1   g543(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n746_), .B(new_n738_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n744_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n745_), .B1(new_n744_), .B2(new_n747_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n731_), .A2(new_n207_), .A3(new_n534_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n667_), .A2(new_n534_), .A3(new_n328_), .A4(new_n704_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(G106gat), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(KEYINPUT114), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n752_), .A3(G106gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(new_n754_), .B2(KEYINPUT114), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n751_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g558(.A(new_n280_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n665_), .A2(new_n760_), .A3(new_n699_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n665_), .A2(KEYINPUT54), .A3(new_n760_), .A4(new_n699_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n305_), .A2(new_n309_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n301_), .A2(new_n297_), .A3(new_n302_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n308_), .C1(new_n295_), .C2(new_n297_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n274_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n256_), .B(new_n257_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n773_), .A2(KEYINPUT55), .A3(new_n247_), .A4(new_n244_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n260_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n244_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n246_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n772_), .B(KEYINPUT56), .C1(new_n779_), .C2(new_n270_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n273_), .A2(new_n310_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n273_), .A2(new_n310_), .A3(KEYINPUT115), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n780_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n779_), .A2(new_n270_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n270_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n772_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n771_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n766_), .B1(new_n792_), .B2(new_n609_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n790_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n270_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n794_), .A2(KEYINPUT116), .A3(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n787_), .A2(KEYINPUT116), .A3(new_n788_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n784_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT115), .B1(new_n273_), .B2(new_n310_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n770_), .B1(new_n796_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(KEYINPUT57), .A3(new_n608_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n273_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT58), .B(new_n804_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n623_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n793_), .A2(new_n803_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n765_), .B1(new_n810_), .B2(new_n328_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n536_), .A2(new_n543_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n578_), .A2(new_n436_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n811_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n310_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT59), .B1(new_n811_), .B2(new_n815_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n810_), .A2(new_n328_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n765_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n814_), .B(KEYINPUT117), .Z(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(KEYINPUT59), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n819_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n824_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n811_), .A2(KEYINPUT118), .A3(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n818_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n310_), .A2(new_n830_), .A3(G113gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n830_), .B2(G113gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n817_), .B1(new_n829_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g632(.A(new_n698_), .ZN(new_n834_));
  OAI21_X1  g633(.A(G120gat), .B1(new_n828_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n836_));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n698_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n816_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(new_n840_), .ZN(G1341gat));
  INV_X1    g640(.A(G127gat), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n328_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n818_), .B(new_n843_), .C1(new_n825_), .C2(new_n827_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n816_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n842_), .B1(new_n845_), .B2(new_n328_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT120), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n844_), .A2(new_n849_), .A3(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(G1342gat));
  OAI21_X1  g650(.A(G134gat), .B1(new_n828_), .B2(new_n665_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n608_), .A2(G134gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n845_), .B2(new_n853_), .ZN(G1343gat));
  NOR3_X1   g653(.A1(new_n690_), .A2(new_n436_), .A3(new_n535_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n822_), .A2(new_n679_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n310_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n384_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n856_), .A2(new_n834_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n385_), .ZN(G1345gat));
  NOR2_X1   g660(.A1(new_n856_), .A2(new_n328_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT61), .B(G155gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  INV_X1    g663(.A(G162gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n856_), .B2(new_n608_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n866_), .A2(KEYINPUT121), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(KEYINPUT121), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n856_), .A2(new_n865_), .A3(new_n665_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(G1347gat));
  NOR3_X1   g669(.A1(new_n679_), .A2(new_n534_), .A3(new_n437_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n822_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT122), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n822_), .A2(new_n874_), .A3(new_n871_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n334_), .A3(new_n310_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G169gat), .B1(new_n872_), .B2(new_n857_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n877_), .B1(new_n879_), .B2(new_n880_), .ZN(G1348gat));
  NAND3_X1  g680(.A1(new_n876_), .A2(new_n335_), .A3(new_n698_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G176gat), .B1(new_n872_), .B2(new_n834_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1349gat));
  NOR3_X1   g683(.A1(new_n872_), .A2(KEYINPUT123), .A3(new_n328_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(G183gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT123), .B1(new_n872_), .B2(new_n328_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n328_), .A2(new_n355_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n886_), .A2(new_n887_), .B1(new_n876_), .B2(new_n888_), .ZN(G1350gat));
  NAND3_X1  g688(.A1(new_n876_), .A2(new_n609_), .A3(new_n356_), .ZN(new_n890_));
  INV_X1    g689(.A(G190gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n665_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1351gat));
  NOR3_X1   g692(.A1(new_n679_), .A2(new_n690_), .A3(new_n573_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n822_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n857_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n450_), .ZN(G1352gat));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n822_), .A2(new_n894_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n834_), .B1(KEYINPUT124), .B2(G204gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n901_), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT125), .B1(new_n895_), .B2(new_n903_), .ZN(new_n904_));
  AND4_X1   g703(.A1(new_n898_), .A2(new_n902_), .A3(new_n453_), .A4(new_n904_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n902_), .A2(new_n904_), .B1(new_n898_), .B2(new_n453_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1353gat));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n908_));
  INV_X1    g707(.A(G211gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n649_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT126), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n899_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n909_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT127), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n912_), .B(new_n914_), .ZN(G1354gat));
  OR3_X1    g714(.A1(new_n895_), .A2(G218gat), .A3(new_n608_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G218gat), .B1(new_n895_), .B2(new_n665_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1355gat));
endmodule


