//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n940_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT3), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT2), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT87), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(KEYINPUT87), .A3(new_n213_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n209_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n207_), .B1(KEYINPUT1), .B2(new_n205_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(KEYINPUT1), .B2(new_n205_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n210_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n212_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n204_), .B1(new_n217_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n216_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n208_), .B1(new_n224_), .B2(new_n214_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n204_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n221_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(KEYINPUT4), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n229_), .B(new_n204_), .C1(new_n217_), .C2(new_n222_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G225gat), .A2(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G1gat), .B(G29gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(G85gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT0), .B(G57gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(new_n237_), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n233_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n234_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n232_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n238_), .B1(new_n243_), .B2(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(G204gat), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT90), .ZN(new_n249_));
  INV_X1    g048(.A(G204gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n250_), .B2(G197gat), .ZN(new_n251_));
  INV_X1    g050(.A(G197gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT21), .B1(new_n248_), .B2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT21), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n246_), .A2(G204gat), .A3(new_n247_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT91), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n252_), .B2(G204gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n260_), .A2(new_n262_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n259_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n264_), .A2(new_n265_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n256_), .A2(new_n259_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n258_), .A2(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G169gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n276_), .B2(new_n272_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n271_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n272_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT83), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(new_n282_), .A3(new_n272_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n272_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n273_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT25), .B(G183gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G190gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G169gat), .ZN(new_n290_));
  INV_X1    g089(.A(G176gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(KEYINPUT24), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT81), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n292_), .A2(KEYINPUT24), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n289_), .A2(new_n299_), .A3(new_n294_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n286_), .A2(new_n296_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n269_), .A2(new_n279_), .A3(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n277_), .A2(new_n297_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n295_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n280_), .A2(KEYINPUT83), .B1(new_n273_), .B2(new_n284_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n278_), .B1(new_n306_), .B2(new_n283_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n271_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n261_), .A2(KEYINPUT91), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n260_), .B(new_n262_), .C1(new_n252_), .C2(G204gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(new_n268_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT21), .B1(new_n310_), .B2(new_n311_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(new_n257_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n302_), .A2(new_n315_), .A3(KEYINPUT20), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n309_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(new_n269_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT20), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n301_), .A2(new_n279_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(new_n314_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n316_), .A2(new_n320_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT95), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n326_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n327_), .B1(new_n326_), .B2(new_n332_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n245_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT92), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n314_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT96), .ZN(new_n338_));
  INV_X1    g137(.A(new_n278_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n308_), .B1(new_n286_), .B2(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n277_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n338_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n305_), .B(KEYINPUT96), .C1(new_n307_), .C2(new_n308_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n312_), .B(KEYINPUT92), .C1(new_n313_), .C2(new_n257_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n337_), .A2(new_n342_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n319_), .B1(new_n345_), .B2(new_n325_), .ZN(new_n346_));
  OAI22_X1  g145(.A1(new_n346_), .A2(KEYINPUT97), .B1(new_n320_), .B2(new_n316_), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n316_), .A2(KEYINPUT97), .A3(new_n320_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n332_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n316_), .A2(new_n320_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n322_), .A2(new_n325_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n331_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n326_), .A2(new_n331_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n223_), .A2(new_n233_), .A3(new_n227_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n239_), .B(new_n356_), .C1(new_n231_), .C2(new_n233_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n244_), .A2(new_n359_), .ZN(new_n360_));
  OAI211_X1 g159(.A(KEYINPUT33), .B(new_n238_), .C1(new_n243_), .C2(new_n240_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OAI22_X1  g161(.A1(new_n335_), .A2(new_n349_), .B1(new_n358_), .B2(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n217_), .A2(new_n222_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n365_), .B(new_n314_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n225_), .B2(new_n221_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n337_), .B2(new_n344_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n368_), .B1(new_n370_), .B2(new_n365_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n225_), .A2(new_n367_), .A3(new_n221_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n373_));
  OR2_X1    g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n373_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G78gat), .B(G106gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT93), .ZN(new_n378_));
  XOR2_X1   g177(.A(G22gat), .B(G50gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n375_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n381_), .B(new_n368_), .C1(new_n370_), .C2(new_n365_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n376_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n376_), .B2(new_n382_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n363_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n352_), .A2(new_n353_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n326_), .A2(new_n331_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n331_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n355_), .A2(KEYINPUT27), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n245_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT99), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n376_), .A2(new_n382_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n380_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n376_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n245_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n355_), .A2(KEYINPUT27), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n347_), .A2(new_n348_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n403_), .B2(new_n331_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT99), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n401_), .A2(new_n404_), .A3(new_n405_), .A4(new_n390_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n386_), .A2(new_n396_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT30), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n324_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n301_), .A2(KEYINPUT30), .A3(new_n279_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(G15gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G71gat), .ZN(new_n415_));
  INV_X1    g214(.A(G99gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT84), .B(G43gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n417_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n419_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT85), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n422_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT85), .B(new_n431_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT86), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n407_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n433_), .A2(new_n245_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n385_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n393_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT64), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT64), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT6), .ZN(new_n448_));
  AND2_X1   g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n446_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G85gat), .ZN(new_n453_));
  INV_X1    g252(.A(G92gat), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n453_), .A2(new_n454_), .A3(KEYINPUT9), .ZN(new_n455_));
  XOR2_X1   g254(.A(G85gat), .B(G92gat), .Z(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(KEYINPUT9), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT10), .B(G99gat), .Z(new_n458_));
  INV_X1    g257(.A(G106gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n452_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT8), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT65), .B1(new_n450_), .B2(new_n451_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n449_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n447_), .A2(KEYINPUT6), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n445_), .A2(KEYINPUT64), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n446_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n463_), .A2(new_n470_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n462_), .B1(new_n475_), .B2(new_n456_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n467_), .A2(new_n469_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n462_), .B(new_n456_), .C1(new_n477_), .C2(new_n473_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n461_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT66), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT15), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT66), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n486_), .B(new_n461_), .C1(new_n476_), .C2(new_n479_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n481_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n489_));
  INV_X1    g288(.A(new_n456_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n473_), .B1(new_n477_), .B2(KEYINPUT65), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n490_), .B1(new_n491_), .B2(new_n470_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n478_), .B1(new_n492_), .B2(new_n462_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(new_n484_), .A3(new_n461_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n488_), .A2(new_n489_), .A3(new_n494_), .A4(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n488_), .A2(new_n489_), .A3(new_n494_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n497_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT35), .B1(new_n488_), .B2(new_n494_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n499_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G190gat), .B(G218gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT69), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT36), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n444_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n488_), .A2(new_n494_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n500_), .B(new_n497_), .C1(new_n510_), .C2(KEYINPUT35), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT71), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n511_), .A2(KEYINPUT72), .A3(new_n499_), .A4(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n511_), .A2(new_n499_), .A3(new_n514_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT72), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(KEYINPUT73), .B(new_n499_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n508_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT73), .B1(new_n511_), .B2(new_n499_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n517_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n525_), .B2(KEYINPUT37), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G57gat), .B(G64gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT11), .ZN(new_n528_));
  XOR2_X1   g327(.A(G71gat), .B(G78gat), .Z(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n528_), .A2(new_n529_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n527_), .A2(KEYINPUT11), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n530_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G1gat), .B(G8gat), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G1gat), .A2(G8gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT14), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n539_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n537_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n544_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(new_n542_), .A3(new_n536_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT75), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n535_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT16), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n535_), .A3(new_n555_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n557_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n561_), .B(new_n562_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n557_), .B2(new_n564_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT76), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT76), .ZN(new_n570_));
  INV_X1    g369(.A(new_n564_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(new_n556_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n565_), .B(new_n570_), .C1(new_n572_), .C2(new_n567_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n526_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n534_), .A2(KEYINPUT12), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n481_), .A2(new_n487_), .A3(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n493_), .A2(new_n461_), .A3(new_n535_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT67), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n480_), .A2(new_n534_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  AOI211_X1 g384(.A(KEYINPUT67), .B(KEYINPUT12), .C1(new_n480_), .C2(new_n534_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n581_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n580_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n535_), .B1(new_n493_), .B2(new_n461_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT5), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n598_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n589_), .A2(new_n593_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT13), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n599_), .A2(KEYINPUT13), .A3(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n545_), .A2(new_n548_), .A3(new_n484_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT78), .Z(new_n610_));
  INV_X1    g409(.A(new_n485_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n608_), .B(new_n610_), .C1(new_n611_), .C2(new_n550_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G113gat), .B(G141gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT79), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G169gat), .B(G197gat), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n614_), .B(new_n615_), .Z(new_n616_));
  AOI21_X1  g415(.A(new_n484_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n617_));
  OAI211_X1 g416(.A(G229gat), .B(G233gat), .C1(new_n607_), .C2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(KEYINPUT77), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(KEYINPUT77), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n612_), .B(new_n616_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT80), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n618_), .B(KEYINPUT77), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT80), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n612_), .A4(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n612_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n616_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n606_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n443_), .A2(new_n576_), .A3(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT100), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n634_), .A2(G1gat), .A3(new_n394_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n407_), .A2(new_n437_), .B1(new_n441_), .B2(new_n439_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n525_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n566_), .A2(new_n568_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n640_), .A3(new_n632_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G1gat), .B1(new_n641_), .B2(new_n394_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n635_), .A2(new_n636_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n637_), .A2(new_n642_), .A3(new_n643_), .ZN(G1324gat));
  INV_X1    g443(.A(new_n393_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G8gat), .B1(new_n641_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n647_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n645_), .A2(G8gat), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n648_), .B(new_n649_), .C1(new_n634_), .C2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g451(.A(new_n437_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n413_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n633_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G15gat), .B1(new_n641_), .B2(new_n437_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT102), .Z(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n657_), .B2(KEYINPUT41), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n658_), .B1(KEYINPUT41), .B2(new_n657_), .ZN(G1326gat));
  OAI21_X1  g458(.A(G22gat), .B1(new_n641_), .B2(new_n385_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n385_), .A2(G22gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n633_), .B2(new_n662_), .ZN(G1327gat));
  NOR3_X1   g462(.A1(new_n638_), .A2(new_n524_), .A3(new_n574_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n632_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n394_), .A2(G29gat), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT105), .Z(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n524_), .A2(new_n444_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n519_), .A2(new_n515_), .A3(new_n509_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n671_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n638_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n526_), .A2(KEYINPUT103), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n516_), .A2(new_n519_), .B1(new_n524_), .B2(new_n444_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n443_), .A2(new_n676_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n675_), .B1(new_n680_), .B2(KEYINPUT43), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n606_), .A2(new_n574_), .A3(new_n631_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n670_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n677_), .B(KEYINPUT103), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n671_), .B1(new_n685_), .B2(new_n443_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n682_), .C1(new_n686_), .C2(new_n675_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n687_), .A3(new_n245_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n684_), .A2(new_n687_), .A3(KEYINPUT104), .A4(new_n245_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G29gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n669_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT106), .B(new_n669_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n665_), .A2(G36gat), .A3(new_n645_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT45), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n684_), .A2(new_n687_), .A3(new_n393_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G36gat), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n699_), .A2(KEYINPUT46), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  XOR2_X1   g505(.A(KEYINPUT107), .B(G43gat), .Z(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n666_), .B2(new_n653_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n684_), .A2(new_n687_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n433_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(G43gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n712_), .B(new_n713_), .Z(G1330gat));
  AOI21_X1  g513(.A(G50gat), .B1(new_n666_), .B2(new_n440_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n440_), .A2(G50gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n709_), .B2(new_n716_), .ZN(G1331gat));
  NOR2_X1   g516(.A1(new_n575_), .A2(new_n630_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n639_), .A2(new_n606_), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G57gat), .B1(new_n719_), .B2(new_n394_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n576_), .A2(new_n606_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(KEYINPUT109), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(KEYINPUT109), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n722_), .A2(new_n443_), .A3(new_n631_), .A4(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT110), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n394_), .A2(G57gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n720_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT111), .B(new_n720_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1332gat));
  OAI21_X1  g530(.A(G64gat), .B1(new_n719_), .B2(new_n645_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT48), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n645_), .A2(G64gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n725_), .B2(new_n734_), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n719_), .B2(new_n437_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT49), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n437_), .A2(G71gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n725_), .B2(new_n738_), .ZN(G1334gat));
  OAI21_X1  g538(.A(G78gat), .B1(new_n719_), .B2(new_n385_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT50), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n385_), .A2(G78gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n725_), .B2(new_n742_), .ZN(G1335gat));
  INV_X1    g542(.A(new_n606_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(new_n630_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n575_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n680_), .A2(KEYINPUT43), .ZN(new_n747_));
  INV_X1    g546(.A(new_n675_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n681_), .A2(KEYINPUT112), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n746_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754_), .B2(new_n394_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n664_), .A2(new_n745_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(new_n453_), .A3(new_n245_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1336gat));
  OAI21_X1  g558(.A(G92gat), .B1(new_n754_), .B2(new_n645_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n454_), .A3(new_n393_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1337gat));
  AOI21_X1  g561(.A(new_n416_), .B1(new_n753_), .B2(new_n653_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n458_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n756_), .A2(new_n764_), .A3(new_n433_), .ZN(new_n765_));
  OR3_X1    g564(.A1(new_n763_), .A2(KEYINPUT51), .A3(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT51), .B1(new_n763_), .B2(new_n765_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1338gat));
  NOR2_X1   g567(.A1(new_n746_), .A2(new_n385_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n459_), .B1(new_n749_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n757_), .A2(new_n459_), .A3(new_n440_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT53), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n772_), .A2(new_n776_), .A3(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1339gat));
  INV_X1    g577(.A(new_n610_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n608_), .B(new_n779_), .C1(new_n611_), .C2(new_n550_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n610_), .B1(new_n607_), .B2(new_n617_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n628_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n601_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT117), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n601_), .A2(new_n783_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n588_), .B1(new_n581_), .B2(new_n587_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n589_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT67), .B1(new_n592_), .B2(KEYINPUT12), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n583_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n792_), .A2(new_n580_), .A3(new_n579_), .A4(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n794_), .A2(new_n790_), .A3(new_n590_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n600_), .B1(new_n791_), .B2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(KEYINPUT56), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n799_), .B(new_n600_), .C1(new_n791_), .C2(new_n796_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n788_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n677_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n788_), .B(KEYINPUT58), .C1(new_n798_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n630_), .A2(new_n601_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n791_), .A2(new_n796_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n598_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n808_), .B1(new_n811_), .B2(new_n800_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n602_), .A2(new_n783_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n806_), .B1(new_n815_), .B2(new_n524_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n790_), .B1(new_n794_), .B2(new_n590_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n794_), .A2(new_n590_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT56), .B(new_n598_), .C1(new_n819_), .C2(new_n795_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n797_), .B2(new_n809_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n813_), .B1(new_n821_), .B2(new_n808_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n822_), .A2(KEYINPUT57), .A3(new_n525_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n805_), .B1(new_n816_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n640_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT57), .B1(new_n822_), .B2(new_n525_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n598_), .B1(new_n819_), .B2(new_n795_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n809_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n807_), .B1(new_n831_), .B2(new_n820_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n806_), .B(new_n524_), .C1(new_n832_), .C2(new_n813_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n828_), .A2(new_n833_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT118), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n826_), .A2(new_n827_), .A3(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n604_), .A2(new_n605_), .A3(new_n718_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n604_), .A2(KEYINPUT114), .A3(new_n605_), .A4(new_n718_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n677_), .A3(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n841_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n836_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n441_), .A2(new_n710_), .A3(new_n245_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n630_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(G113gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(KEYINPUT119), .A3(new_n851_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n824_), .A2(new_n856_), .A3(new_n575_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT120), .B1(new_n834_), .B2(new_n574_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n846_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n848_), .A2(KEYINPUT59), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n848_), .B1(new_n836_), .B2(new_n846_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n631_), .A2(new_n851_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n854_), .A2(new_n855_), .B1(new_n865_), .B2(new_n866_), .ZN(G1340gat));
  OAI21_X1  g666(.A(G120gat), .B1(new_n864_), .B2(new_n744_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n862_), .ZN(new_n869_));
  INV_X1    g668(.A(G120gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n744_), .B2(KEYINPUT60), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(KEYINPUT60), .B2(new_n870_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n869_), .B2(new_n872_), .ZN(G1341gat));
  OAI21_X1  g672(.A(G127gat), .B1(new_n864_), .B2(new_n827_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n575_), .A2(G127gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n869_), .B2(new_n875_), .ZN(G1342gat));
  AOI21_X1  g675(.A(G134gat), .B1(new_n862_), .B2(new_n525_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT121), .B(G134gat), .Z(new_n878_));
  NAND2_X1  g677(.A1(new_n526_), .A2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT122), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n877_), .B1(new_n865_), .B2(new_n880_), .ZN(G1343gat));
  NOR4_X1   g680(.A1(new_n653_), .A2(new_n394_), .A3(new_n385_), .A4(new_n393_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n847_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n631_), .ZN(new_n884_));
  INV_X1    g683(.A(G141gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1344gat));
  NOR2_X1   g685(.A1(new_n883_), .A2(new_n744_), .ZN(new_n887_));
  INV_X1    g686(.A(G148gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1345gat));
  NOR2_X1   g688(.A1(new_n883_), .A2(new_n575_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT61), .B(G155gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  AND2_X1   g691(.A1(new_n847_), .A2(new_n882_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G162gat), .B1(new_n893_), .B2(new_n525_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n685_), .A2(G162gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n893_), .B2(new_n895_), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n645_), .A2(new_n245_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n653_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n440_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n630_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n841_), .A2(new_n845_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n824_), .A2(new_n575_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(KEYINPUT120), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n900_), .B1(new_n904_), .B2(new_n857_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n905_), .C2(new_n290_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  INV_X1    g706(.A(new_n900_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n290_), .B1(new_n859_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n907_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n290_), .A2(KEYINPUT62), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT123), .B1(new_n905_), .B2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n859_), .A2(new_n908_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n916_), .A3(new_n912_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n906_), .A2(new_n911_), .A3(new_n914_), .A4(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT22), .B(G169gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n905_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1348gat));
  NAND2_X1  g720(.A1(new_n847_), .A2(new_n385_), .ZN(new_n922_));
  NOR4_X1   g721(.A1(new_n922_), .A2(new_n291_), .A3(new_n744_), .A4(new_n898_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n859_), .A2(new_n606_), .A3(new_n899_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n291_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n924_), .A2(KEYINPUT125), .A3(new_n291_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n923_), .B1(new_n927_), .B2(new_n928_), .ZN(G1349gat));
  AND2_X1   g728(.A1(new_n859_), .A2(new_n899_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n827_), .A2(new_n287_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(KEYINPUT126), .A3(new_n931_), .ZN(new_n935_));
  INV_X1    g734(.A(G183gat), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n653_), .A2(new_n574_), .A3(new_n897_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n922_), .B2(new_n937_), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n934_), .A2(new_n935_), .A3(new_n938_), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n930_), .A2(new_n525_), .A3(new_n288_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n930_), .A2(new_n526_), .ZN(new_n941_));
  INV_X1    g740(.A(G190gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(G1351gat));
  NAND3_X1  g742(.A1(new_n437_), .A2(new_n401_), .A3(new_n393_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n944_), .B1(new_n836_), .B2(new_n846_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n630_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n606_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g748(.A(KEYINPUT63), .B(G211gat), .C1(new_n945_), .C2(new_n640_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n945_), .A2(new_n640_), .ZN(new_n951_));
  XOR2_X1   g750(.A(KEYINPUT63), .B(G211gat), .Z(new_n952_));
  AOI21_X1  g751(.A(new_n950_), .B1(new_n951_), .B2(new_n952_), .ZN(G1354gat));
  AOI21_X1  g752(.A(G218gat), .B1(new_n945_), .B2(new_n525_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n526_), .A2(G218gat), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(KEYINPUT127), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n954_), .B1(new_n945_), .B2(new_n956_), .ZN(G1355gat));
endmodule


