//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G85gat), .B(G92gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT6), .ZN(new_n206_));
  OR4_X1    g005(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT7), .ZN(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT66), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n207_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n214_), .B(KEYINPUT65), .Z(new_n215_));
  OAI21_X1  g014(.A(new_n204_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n204_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G85gat), .B(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(KEYINPUT9), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n222_), .A3(KEYINPUT64), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT10), .B(G99gat), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n210_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n225_), .A2(new_n206_), .A3(new_n226_), .A4(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n217_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G57gat), .B(G64gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT67), .ZN(new_n233_));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(KEYINPUT11), .B2(new_n231_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n233_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n230_), .A2(new_n236_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n203_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n240_), .A2(KEYINPUT68), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n236_), .B(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n229_), .A2(KEYINPUT69), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n229_), .A2(KEYINPUT69), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n217_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n247_), .A2(new_n237_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n239_), .A2(KEYINPUT12), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n202_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(KEYINPUT68), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n241_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G120gat), .B(G148gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT5), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G176gat), .B(G204gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n254_), .B(new_n255_), .Z(new_n256_));
  NOR2_X1   g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT72), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n256_), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT71), .Z(new_n260_));
  INV_X1    g059(.A(KEYINPUT13), .ZN(new_n261_));
  OR3_X1    g060(.A1(new_n258_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n261_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G1gat), .B(G8gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT78), .ZN(new_n269_));
  INV_X1    g068(.A(G15gat), .ZN(new_n270_));
  INV_X1    g069(.A(G22gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G15gat), .A2(G22gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G1gat), .A2(G8gat), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n272_), .A2(new_n273_), .B1(KEYINPUT14), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n269_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G29gat), .B(G36gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT74), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G43gat), .B(G50gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(KEYINPUT15), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n283_), .B2(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G229gat), .A2(G233gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(KEYINPUT81), .Z(new_n286_));
  XOR2_X1   g085(.A(new_n281_), .B(new_n276_), .Z(new_n287_));
  INV_X1    g086(.A(new_n285_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n284_), .A2(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G113gat), .B(G141gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT82), .ZN(new_n291_));
  XOR2_X1   g090(.A(G169gat), .B(G197gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT83), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n289_), .A2(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n230_), .A2(new_n281_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G232gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT34), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(KEYINPUT35), .B2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n246_), .B2(new_n283_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(KEYINPUT35), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G190gat), .B(G218gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT75), .ZN(new_n307_));
  XOR2_X1   g106(.A(G134gat), .B(G162gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  OR3_X1    g109(.A1(new_n305_), .A2(KEYINPUT36), .A3(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n309_), .B(KEYINPUT36), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n305_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT37), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n315_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT77), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n317_), .A2(new_n318_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n314_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n317_), .A2(new_n318_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n314_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G231gat), .A2(G233gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT79), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n236_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(new_n277_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G155gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT16), .ZN(new_n333_));
  XOR2_X1   g132(.A(G183gat), .B(G211gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(KEYINPUT70), .A3(KEYINPUT17), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n331_), .A2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(KEYINPUT17), .B2(new_n336_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n330_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n326_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT80), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n326_), .A2(new_n344_), .A3(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n267_), .A2(new_n298_), .A3(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(KEYINPUT86), .A2(G183gat), .A3(G190gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT86), .B1(G183gat), .B2(G190gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT23), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT88), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n350_), .A2(new_n357_), .A3(new_n351_), .A4(new_n354_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n359_));
  AOI21_X1  g158(.A(G176gat), .B1(new_n359_), .B2(KEYINPUT22), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G169gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n356_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n353_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n352_), .A2(KEYINPUT23), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OR3_X1    g164(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n366_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT26), .B(G190gat), .ZN(new_n372_));
  INV_X1    g171(.A(G183gat), .ZN(new_n373_));
  OR2_X1    g172(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n374_));
  NAND2_X1  g173(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n372_), .B1(new_n376_), .B2(KEYINPUT85), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378_));
  INV_X1    g177(.A(new_n375_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n380_));
  OAI21_X1  g179(.A(G183gat), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n373_), .A2(KEYINPUT25), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n378_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n365_), .B(new_n371_), .C1(new_n377_), .C2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n362_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G71gat), .B(G99gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(G43gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n385_), .B(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G127gat), .B(G134gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(G113gat), .B(G120gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n388_), .B(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(new_n270_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT30), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT31), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n392_), .B(new_n396_), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT89), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(KEYINPUT1), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n402_), .B2(KEYINPUT1), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT91), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n404_), .B2(new_n403_), .ZN(new_n406_));
  AND3_X1   g205(.A1(KEYINPUT90), .A2(G141gat), .A3(G148gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G141gat), .ZN(new_n410_));
  INV_X1    g209(.A(G148gat), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT92), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT92), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n420_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT2), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n400_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(new_n402_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n425_), .A2(KEYINPUT93), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT93), .B1(new_n425_), .B2(new_n427_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n413_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT94), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT94), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n413_), .B(new_n432_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435_));
  OR3_X1    g234(.A1(new_n434_), .A2(KEYINPUT96), .A3(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(G228gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT21), .ZN(new_n439_));
  INV_X1    g238(.A(G204gat), .ZN(new_n440_));
  OR2_X1    g239(.A1(KEYINPUT97), .A2(G197gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(KEYINPUT97), .A2(G197gat), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G197gat), .A2(G204gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n439_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G211gat), .B(G218gat), .Z(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n439_), .B1(G197gat), .B2(G204gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n446_), .A2(KEYINPUT21), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n443_), .A2(new_n444_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n445_), .A2(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT96), .B1(new_n434_), .B2(new_n435_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n436_), .A2(new_n438_), .A3(new_n453_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n430_), .A2(KEYINPUT29), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n438_), .B1(new_n456_), .B2(new_n453_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G22gat), .B(G50gat), .Z(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n463_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n464_));
  AOI211_X1 g263(.A(KEYINPUT29), .B(new_n462_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n461_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n464_), .A2(new_n465_), .A3(new_n461_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G78gat), .B(G106gat), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(KEYINPUT98), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n464_), .A2(new_n465_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n461_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n471_), .B1(new_n474_), .B2(new_n466_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n460_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n469_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n477_), .A3(new_n466_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n467_), .A2(new_n468_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n459_), .B(new_n478_), .C1(new_n479_), .C2(new_n471_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G29gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(G85gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT0), .B(G57gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  NAND3_X1  g284(.A1(new_n431_), .A2(new_n433_), .A3(new_n391_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n430_), .A2(new_n391_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n487_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G225gat), .A2(G233gat), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n489_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n486_), .A2(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n492_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n485_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(KEYINPUT4), .ZN(new_n498_));
  INV_X1    g297(.A(new_n492_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n488_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n485_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n495_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(KEYINPUT109), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT109), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n500_), .A2(new_n504_), .A3(new_n501_), .A4(new_n495_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT18), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G64gat), .B(G92gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT32), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT101), .ZN(new_n511_));
  INV_X1    g310(.A(G169gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT22), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT22), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(G169gat), .ZN(new_n515_));
  INV_X1    g314(.A(G176gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n513_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n367_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT99), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n352_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(KEYINPUT86), .A2(G183gat), .A3(G190gat), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT23), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n364_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n351_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT99), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n517_), .A2(new_n526_), .A3(new_n367_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n519_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT25), .B(G183gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n372_), .A2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n371_), .A2(new_n354_), .A3(new_n350_), .A4(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n511_), .B1(new_n532_), .B2(new_n453_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n528_), .A2(new_n531_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(KEYINPUT101), .A3(new_n452_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n385_), .A2(new_n453_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G226gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT19), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .A4(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT20), .B1(new_n385_), .B2(new_n453_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT100), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n534_), .B2(new_n452_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n453_), .A2(new_n532_), .A3(KEYINPUT100), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n542_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n538_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n541_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT106), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n510_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT32), .B(new_n509_), .C1(new_n548_), .C2(KEYINPUT106), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n360_), .B(new_n512_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(KEYINPUT88), .B2(new_n355_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n382_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT85), .B1(new_n376_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n381_), .A2(new_n378_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n372_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n370_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n553_), .A2(new_n358_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n539_), .B1(new_n559_), .B2(new_n452_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n453_), .A2(new_n532_), .A3(KEYINPUT100), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT100), .B1(new_n453_), .B2(new_n532_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n560_), .B(new_n547_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT108), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n544_), .A2(new_n545_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT108), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n547_), .A4(new_n560_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT107), .B(KEYINPUT20), .Z(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n534_), .B2(new_n452_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n547_), .B1(new_n569_), .B2(new_n536_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(new_n567_), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n550_), .B1(new_n551_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n503_), .A2(new_n505_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT110), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n503_), .A2(KEYINPUT110), .A3(new_n505_), .A4(new_n573_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n501_), .B1(new_n500_), .B2(new_n495_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(KEYINPUT104), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT104), .ZN(new_n582_));
  AOI211_X1 g381(.A(new_n582_), .B(new_n501_), .C1(new_n500_), .C2(new_n495_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT105), .B1(new_n581_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n497_), .A2(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(KEYINPUT104), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT105), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .A4(new_n579_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT33), .B(new_n485_), .C1(new_n493_), .C2(new_n496_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n509_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n548_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT103), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT103), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n548_), .A2(new_n593_), .A3(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n492_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n596_), .B(new_n501_), .C1(new_n494_), .C2(new_n492_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n509_), .B(new_n541_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT102), .ZN(new_n599_));
  AND4_X1   g398(.A1(new_n589_), .A2(new_n595_), .A3(new_n597_), .A4(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n584_), .A2(new_n588_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n481_), .B1(new_n578_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n503_), .A2(new_n505_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n481_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(new_n599_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT27), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n572_), .A2(KEYINPUT111), .A3(new_n590_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n598_), .A2(KEYINPUT27), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT111), .B1(new_n572_), .B2(new_n590_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n611_), .A2(KEYINPUT112), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT112), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n570_), .B1(new_n563_), .B2(KEYINPUT108), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n509_), .B1(new_n615_), .B2(new_n567_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n609_), .B1(new_n616_), .B2(KEYINPUT111), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n572_), .A2(new_n590_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT111), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n614_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n607_), .B1(new_n613_), .B2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n604_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(KEYINPUT113), .B(new_n399_), .C1(new_n602_), .C2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT113), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n601_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n481_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n628_), .B2(new_n398_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n624_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n622_), .A2(new_n481_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n603_), .A2(new_n397_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n347_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n603_), .A2(G1gat), .ZN(new_n637_));
  OR3_X1    g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n298_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n264_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n341_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n324_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n634_), .A3(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n603_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n636_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n638_), .A2(new_n644_), .A3(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n622_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n648_), .A2(new_n649_), .A3(G8gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n648_), .B2(G8gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n622_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(G8gat), .ZN(new_n653_));
  OAI22_X1  g452(.A1(new_n650_), .A2(new_n651_), .B1(new_n635_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT114), .B(KEYINPUT40), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n654_), .B(new_n656_), .ZN(G1325gat));
  INV_X1    g456(.A(new_n635_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n270_), .A3(new_n398_), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT115), .B(KEYINPUT41), .Z(new_n660_));
  NAND2_X1  g459(.A1(new_n647_), .A2(new_n398_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(G15gat), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n661_), .A2(G15gat), .A3(new_n660_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(G1326gat));
  NAND3_X1  g463(.A1(new_n658_), .A2(new_n271_), .A3(new_n481_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT116), .B(KEYINPUT42), .Z(new_n666_));
  NAND2_X1  g465(.A1(new_n647_), .A2(new_n481_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(G22gat), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(G22gat), .A3(new_n666_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1327gat));
  NOR2_X1   g469(.A1(new_n314_), .A2(new_n341_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n640_), .A2(new_n634_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n603_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G29gat), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n326_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(KEYINPUT117), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT117), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n624_), .A2(new_n629_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n678_), .B(KEYINPUT43), .C1(new_n679_), .C2(new_n326_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n640_), .A2(new_n641_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT44), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  AOI211_X1 g484(.A(new_n685_), .B(new_n682_), .C1(new_n677_), .C2(new_n680_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n673_), .A2(G29gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n674_), .B1(new_n687_), .B2(new_n688_), .ZN(G1328gat));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  INV_X1    g489(.A(G36gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n687_), .B2(new_n622_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n622_), .B(KEYINPUT118), .Z(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n672_), .A2(new_n691_), .A3(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT45), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n690_), .B1(new_n692_), .B2(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n684_), .A2(new_n686_), .A3(new_n652_), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT46), .B(new_n696_), .C1(new_n699_), .C2(new_n691_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n681_), .A2(new_n683_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n685_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n683_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n397_), .A2(G43gat), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G43gat), .B1(new_n672_), .B2(new_n398_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT47), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n687_), .B2(new_n705_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(G1330gat));
  INV_X1    g511(.A(G50gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n672_), .A2(new_n713_), .A3(new_n481_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n703_), .A2(new_n481_), .A3(new_n704_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT119), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(G50gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n715_), .B2(G50gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1331gat));
  NOR2_X1   g518(.A1(new_n679_), .A2(new_n298_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n266_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n642_), .ZN(new_n722_));
  INV_X1    g521(.A(G57gat), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n603_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n346_), .A2(new_n264_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT120), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n720_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT121), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT121), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(new_n730_), .A3(new_n720_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n729_), .A2(new_n673_), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n724_), .B1(new_n732_), .B2(new_n723_), .ZN(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n722_), .B2(new_n693_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n693_), .A2(G64gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n728_), .B2(new_n736_), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n722_), .B2(new_n399_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT49), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n399_), .A2(G71gat), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT122), .Z(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n728_), .B2(new_n741_), .ZN(G1334gat));
  NAND3_X1  g541(.A1(new_n721_), .A2(new_n642_), .A3(new_n481_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(G78gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(G78gat), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n627_), .A2(G78gat), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n745_), .A2(new_n746_), .B1(new_n728_), .B2(new_n747_), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n721_), .A2(new_n671_), .ZN(new_n749_));
  OR3_X1    g548(.A1(new_n749_), .A2(G85gat), .A3(new_n603_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n264_), .A2(new_n641_), .A3(new_n639_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n677_), .B2(new_n680_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753_), .B2(new_n603_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n750_), .A2(new_n754_), .ZN(G1336gat));
  INV_X1    g554(.A(new_n749_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n221_), .A3(new_n622_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G92gat), .B1(new_n753_), .B2(new_n693_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1337gat));
  AND4_X1   g558(.A1(new_n227_), .A2(new_n721_), .A3(new_n397_), .A4(new_n671_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n209_), .B1(new_n752_), .B2(new_n398_), .ZN(new_n761_));
  OAI22_X1  g560(.A1(new_n760_), .A2(new_n761_), .B1(KEYINPUT123), .B2(KEYINPUT51), .ZN(new_n762_));
  NAND2_X1  g561(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n756_), .A2(new_n210_), .A3(new_n481_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT124), .B(KEYINPUT52), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n752_), .A2(new_n481_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G106gat), .ZN(new_n768_));
  INV_X1    g567(.A(new_n766_), .ZN(new_n769_));
  AOI211_X1 g568(.A(new_n210_), .B(new_n769_), .C1(new_n752_), .C2(new_n481_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n765_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n765_), .B(new_n773_), .C1(new_n768_), .C2(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  NAND3_X1  g574(.A1(new_n262_), .A2(new_n639_), .A3(new_n263_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n342_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n342_), .A2(new_n776_), .A3(KEYINPUT54), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n286_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n284_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n293_), .B1(new_n287_), .B2(new_n286_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n295_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n258_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n248_), .A2(new_n249_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n203_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(new_n250_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n256_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(KEYINPUT56), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n791_), .A2(new_n795_), .A3(new_n792_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n787_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n786_), .B1(new_n797_), .B2(new_n639_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n314_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(KEYINPUT57), .A3(new_n314_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n787_), .B(new_n785_), .C1(new_n794_), .C2(new_n796_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n322_), .A2(new_n325_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT125), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n803_), .A2(new_n804_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n807_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n801_), .B(new_n802_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n781_), .B1(new_n812_), .B2(new_n641_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n631_), .A2(new_n673_), .A3(new_n397_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n298_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n641_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n781_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n821_), .A2(KEYINPUT126), .ZN(new_n822_));
  INV_X1    g621(.A(new_n814_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(KEYINPUT126), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT126), .B(new_n821_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n639_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n817_), .B1(new_n827_), .B2(new_n816_), .ZN(G1340gat));
  INV_X1    g627(.A(KEYINPUT60), .ZN(new_n829_));
  AOI21_X1  g628(.A(G120gat), .B1(new_n264_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n829_), .B2(G120gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n815_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n267_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n833_));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(G1341gat));
  INV_X1    g634(.A(G127gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n815_), .A2(new_n836_), .A3(new_n341_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n641_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n836_), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n815_), .A2(new_n840_), .A3(new_n324_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n326_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n840_), .ZN(G1343gat));
  NOR2_X1   g642(.A1(new_n627_), .A2(new_n398_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n694_), .A2(new_n603_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n820_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n410_), .A3(new_n298_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G141gat), .B1(new_n846_), .B2(new_n639_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1344gat));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n411_), .A3(new_n266_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G148gat), .B1(new_n846_), .B2(new_n267_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1345gat));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  OR3_X1    g653(.A1(new_n846_), .A2(new_n641_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n846_), .B2(new_n641_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1346gat));
  OAI21_X1  g656(.A(G162gat), .B1(new_n846_), .B2(new_n326_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n314_), .A2(G162gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n846_), .B2(new_n859_), .ZN(G1347gat));
  NOR4_X1   g659(.A1(new_n693_), .A2(new_n673_), .A3(new_n481_), .A4(new_n399_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n820_), .A2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G169gat), .B1(new_n862_), .B2(new_n639_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT62), .B(G169gat), .C1(new_n862_), .C2(new_n639_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n862_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n867_), .A2(new_n298_), .A3(new_n513_), .A4(new_n515_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n866_), .A3(new_n868_), .ZN(G1348gat));
  OAI21_X1  g668(.A(G176gat), .B1(new_n862_), .B2(new_n267_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n264_), .A2(new_n516_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n862_), .B2(new_n871_), .ZN(G1349gat));
  NAND3_X1  g671(.A1(new_n867_), .A2(new_n341_), .A3(new_n529_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G183gat), .B1(new_n862_), .B2(new_n641_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1350gat));
  OAI21_X1  g674(.A(G190gat), .B1(new_n862_), .B2(new_n326_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n324_), .A2(new_n372_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n862_), .B2(new_n877_), .ZN(G1351gat));
  NOR2_X1   g677(.A1(new_n693_), .A2(new_n673_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n820_), .A2(new_n844_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G197gat), .B1(new_n881_), .B2(new_n298_), .ZN(new_n882_));
  INV_X1    g681(.A(G197gat), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n880_), .A2(new_n883_), .A3(new_n639_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1352gat));
  NAND3_X1  g684(.A1(new_n881_), .A2(new_n440_), .A3(new_n266_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G204gat), .B1(new_n880_), .B2(new_n267_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1353gat));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n341_), .A2(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT127), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n881_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n893_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n880_), .A2(new_n889_), .A3(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1354gat));
  OAI21_X1  g696(.A(G218gat), .B1(new_n880_), .B2(new_n326_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n314_), .A2(G218gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n880_), .B2(new_n899_), .ZN(G1355gat));
endmodule


