//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_;
  XNOR2_X1  g000(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT81), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT81), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G169gat), .A3(G176gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT82), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT23), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n215_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n210_), .B(new_n214_), .C1(new_n219_), .C2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(KEYINPUT25), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G190gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n226_), .B(new_n228_), .C1(KEYINPUT80), .C2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n225_), .A2(KEYINPUT25), .ZN(new_n232_));
  INV_X1    g031(.A(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT26), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(KEYINPUT26), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n232_), .B(new_n234_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n231_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n221_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n220_), .A2(KEYINPUT23), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243_));
  OAI21_X1  g042(.A(G169gat), .B1(new_n243_), .B2(KEYINPUT83), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n212_), .A2(KEYINPUT22), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n244_), .B(new_n213_), .C1(KEYINPUT83), .C2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n207_), .A2(new_n209_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  OAI22_X1  g048(.A1(new_n223_), .A2(new_n238_), .B1(new_n242_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n251_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G15gat), .B(G43gat), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n254_), .A2(new_n255_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n203_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n202_), .A3(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G227gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(G71gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n259_), .A2(new_n261_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G113gat), .B(G120gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(G127gat), .B(G134gat), .Z(new_n269_));
  INV_X1    g068(.A(KEYINPUT87), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G127gat), .B(G134gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT87), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n268_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n273_), .A3(new_n268_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT86), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n278_), .B2(new_n277_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G99gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n266_), .A2(new_n267_), .A3(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n282_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G226gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n239_), .A2(new_n241_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n206_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n214_), .B1(new_n290_), .B2(new_n204_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT25), .B(G183gat), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n230_), .A2(new_n234_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n240_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT22), .B(G169gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n247_), .B1(new_n213_), .B2(new_n297_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n289_), .A2(new_n294_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G197gat), .B(G204gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301_));
  OAI211_X1 g100(.A(KEYINPUT21), .B(new_n300_), .C1(new_n301_), .C2(KEYINPUT90), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT21), .ZN(new_n303_));
  INV_X1    g102(.A(G218gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G211gat), .ZN(new_n305_));
  INV_X1    g104(.A(G211gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G218gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT90), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n303_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(G197gat), .A2(G204gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G197gat), .A2(G204gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(new_n301_), .B2(KEYINPUT21), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n302_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT20), .B1(new_n299_), .B2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n250_), .A2(new_n315_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n288_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT20), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n299_), .B2(new_n316_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n288_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n250_), .A2(new_n315_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n319_), .A2(KEYINPUT93), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT93), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n326_), .B(new_n288_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT18), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n317_), .A2(new_n318_), .A3(new_n288_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n322_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n332_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n334_), .A2(KEYINPUT27), .A3(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G155gat), .B(G162gat), .Z(new_n340_));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(G141gat), .ZN(new_n344_));
  INV_X1    g143(.A(G148gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n342_), .A2(new_n343_), .A3(new_n346_), .A4(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT88), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n343_), .A2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n350_), .B(new_n351_), .C1(new_n353_), .C2(KEYINPUT2), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n353_), .A2(KEYINPUT2), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n340_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n348_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT29), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n315_), .ZN(new_n359_));
  AND2_X1   g158(.A1(G228gat), .A2(G233gat), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n360_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT91), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n367_));
  OR3_X1    g166(.A1(new_n357_), .A2(KEYINPUT29), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n357_), .B2(KEYINPUT29), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G22gat), .B(G50gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n366_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n361_), .A2(new_n362_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n363_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n365_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n366_), .A2(new_n372_), .A3(new_n375_), .A4(new_n365_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT96), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n357_), .A2(new_n276_), .A3(new_n275_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n271_), .A2(new_n273_), .A3(new_n268_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n356_), .B(new_n348_), .C1(new_n383_), .C2(new_n274_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n384_), .A3(KEYINPUT4), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n357_), .A2(new_n275_), .A3(new_n386_), .A4(new_n276_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n381_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n380_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391_));
  INV_X1    g190(.A(G85gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n390_), .A2(new_n395_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n377_), .A2(new_n378_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n325_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n334_), .A2(KEYINPUT94), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n325_), .A2(new_n402_), .A3(new_n327_), .A4(new_n332_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT98), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n400_), .A2(KEYINPUT98), .A3(new_n401_), .A4(new_n403_), .ZN(new_n407_));
  AOI211_X1 g206(.A(new_n339_), .B(new_n398_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n377_), .A2(new_n378_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n325_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n332_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n402_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n403_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n411_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n400_), .A2(KEYINPUT95), .A3(new_n403_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n385_), .A2(new_n387_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n395_), .B1(new_n418_), .B2(new_n381_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n382_), .A2(new_n384_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n381_), .B1(new_n420_), .B2(KEYINPUT97), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(KEYINPUT97), .B2(new_n420_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n424_), .B(new_n395_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n423_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n416_), .A2(new_n417_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n397_), .A2(new_n396_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT32), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n328_), .B1(new_n432_), .B2(new_n332_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n337_), .A2(KEYINPUT32), .A3(new_n333_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n410_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n285_), .B1(new_n408_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT99), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n285_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n431_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n339_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n440_), .A2(new_n409_), .A3(new_n441_), .A4(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(KEYINPUT99), .B(new_n285_), .C1(new_n408_), .C2(new_n436_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n439_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G15gat), .B(G22gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT74), .ZN(new_n447_));
  INV_X1    g246(.A(G1gat), .ZN(new_n448_));
  INV_X1    g247(.A(G8gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT14), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n447_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT75), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n453_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT75), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n451_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G1gat), .B(G8gat), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n454_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G43gat), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT15), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n462_), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT78), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G229gat), .A2(G233gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n461_), .A2(new_n462_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n471_), .B2(new_n465_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n465_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n468_), .A2(new_n472_), .B1(new_n473_), .B2(new_n470_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G113gat), .B(G141gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G169gat), .B(G197gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n474_), .B(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n445_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(G92gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n392_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G85gat), .A2(G92gat), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT6), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(G99gat), .A3(G106gat), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n489_));
  INV_X1    g288(.A(G99gat), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n483_), .B1(new_n488_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT66), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n485_), .A2(new_n487_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(new_n493_), .A3(new_n492_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n483_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n496_), .A2(KEYINPUT8), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT65), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n481_), .A2(new_n502_), .A3(KEYINPUT9), .A4(new_n482_), .ZN(new_n503_));
  OR2_X1    g302(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n491_), .A3(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n503_), .A2(new_n497_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT9), .ZN(new_n508_));
  INV_X1    g307(.A(new_n482_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n508_), .B(new_n481_), .C1(new_n509_), .C2(KEYINPUT65), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n496_), .B2(KEYINPUT8), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n501_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n465_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G232gat), .A2(G233gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT34), .Z(new_n516_));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT71), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n499_), .B1(new_n498_), .B2(new_n483_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n523_), .A2(new_n524_), .B1(new_n510_), .B2(new_n507_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n496_), .A2(KEYINPUT8), .A3(new_n500_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT67), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n466_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT67), .B1(new_n501_), .B2(new_n512_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n466_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT70), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n514_), .A2(KEYINPUT72), .A3(new_n519_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n522_), .A2(new_n532_), .A3(new_n536_), .A4(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n516_), .A2(new_n517_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n520_), .A2(new_n539_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n535_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT73), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G134gat), .B(G162gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT36), .Z(new_n548_));
  NAND3_X1  g347(.A1(new_n543_), .A2(new_n544_), .A3(new_n548_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n538_), .A2(new_n539_), .B1(new_n535_), .B2(new_n541_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n548_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT73), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n547_), .A2(KEYINPUT36), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT37), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n543_), .A2(new_n548_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n555_), .A2(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n562_));
  XOR2_X1   g361(.A(G71gat), .B(G78gat), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(KEYINPUT12), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n533_), .A2(new_n534_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n565_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n501_), .B2(new_n512_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n533_), .A2(KEYINPUT68), .A3(new_n534_), .A4(new_n567_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT64), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n513_), .B2(new_n571_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n570_), .A2(new_n575_), .A3(new_n576_), .A4(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n513_), .A2(new_n571_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n573_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n578_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G120gat), .B(G148gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n589_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n580_), .A2(new_n583_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(KEYINPUT13), .A3(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n471_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n571_), .B(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n471_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT77), .B1(new_n603_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT17), .B1(new_n602_), .B2(new_n605_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n615_), .B1(new_n616_), .B2(new_n613_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n608_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n559_), .A2(new_n598_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n479_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(new_n448_), .A3(new_n431_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n478_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n597_), .A2(new_n629_), .A3(new_n620_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n445_), .A2(new_n555_), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n441_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n627_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n628_), .A2(new_n632_), .A3(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n442_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n625_), .A2(new_n449_), .A3(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n631_), .A2(new_n442_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n449_), .B1(new_n637_), .B2(KEYINPUT100), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n631_), .B2(new_n442_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n639_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n636_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT40), .B(new_n636_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n631_), .B2(new_n285_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT41), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n624_), .A2(G15gat), .A3(new_n285_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1326gat));
  OAI21_X1  g451(.A(G22gat), .B1(new_n631_), .B2(new_n409_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT42), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n409_), .A2(G22gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n624_), .B2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(new_n555_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n620_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n597_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n479_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G29gat), .B1(new_n661_), .B2(new_n431_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n559_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n444_), .A2(new_n443_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n406_), .A2(new_n407_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n339_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n398_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n400_), .A2(new_n403_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n428_), .B1(new_n670_), .B2(new_n411_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n671_), .B2(new_n417_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n410_), .B2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT99), .B1(new_n673_), .B2(new_n285_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n663_), .B1(new_n664_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT43), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n677_), .B(new_n663_), .C1(new_n664_), .C2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n598_), .A2(new_n478_), .A3(new_n620_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT102), .Z(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT44), .B1(new_n679_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n684_), .B(new_n681_), .C1(new_n676_), .C2(new_n678_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n431_), .A2(G29gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n662_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  INV_X1    g488(.A(G36gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n686_), .B2(new_n635_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n635_), .A2(new_n690_), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n660_), .A2(KEYINPUT45), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT45), .B1(new_n660_), .B2(new_n692_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n689_), .B1(new_n691_), .B2(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n683_), .A2(new_n685_), .A3(new_n442_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT46), .B(new_n695_), .C1(new_n698_), .C2(new_n690_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1329gat));
  INV_X1    g499(.A(G43gat), .ZN(new_n701_));
  NOR4_X1   g500(.A1(new_n683_), .A2(new_n685_), .A3(new_n701_), .A4(new_n285_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G43gat), .B1(new_n661_), .B2(new_n440_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT47), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n285_), .A2(new_n701_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n686_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n704_), .A2(new_n708_), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n661_), .B2(new_n410_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n410_), .A2(G50gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n686_), .B2(new_n711_), .ZN(G1331gat));
  AND2_X1   g511(.A1(new_n445_), .A2(new_n629_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n559_), .A2(new_n597_), .A3(new_n621_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT103), .Z(new_n715_));
  AND2_X1   g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(G57gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n431_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n445_), .A2(new_n555_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n598_), .A2(new_n478_), .A3(new_n620_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n441_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT104), .Z(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n716_), .A2(new_n725_), .A3(new_n635_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n721_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n727_), .B2(new_n635_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT105), .B(KEYINPUT48), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n729_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n730_), .B2(new_n731_), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n721_), .B2(new_n285_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT49), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n716_), .A2(new_n263_), .A3(new_n440_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1334gat));
  OAI21_X1  g535(.A(G78gat), .B1(new_n721_), .B2(new_n409_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT50), .ZN(new_n738_));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n716_), .A2(new_n739_), .A3(new_n410_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n658_), .A2(new_n598_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n713_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n392_), .A3(new_n431_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n598_), .A2(new_n478_), .A3(new_n621_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n678_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n677_), .B1(new_n445_), .B2(new_n663_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT106), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n679_), .A2(new_n751_), .A3(new_n746_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n441_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n745_), .B1(new_n753_), .B2(new_n392_), .ZN(G1336gat));
  OAI21_X1  g553(.A(new_n480_), .B1(new_n743_), .B2(new_n442_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT107), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n750_), .A2(new_n752_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n442_), .A2(new_n480_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(G1337gat));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n440_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n743_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n743_), .B2(new_n761_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n285_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n490_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT51), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n764_), .B(new_n768_), .C1(new_n765_), .C2(new_n490_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n744_), .A2(new_n491_), .A3(new_n410_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n679_), .A2(new_n410_), .A3(new_n746_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n773_), .A3(G106gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(G106gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n771_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  NOR2_X1   g579(.A1(new_n635_), .A2(new_n410_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n285_), .A2(new_n441_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n478_), .A2(new_n592_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT68), .B1(new_n530_), .B2(new_n567_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n576_), .A2(new_n575_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(KEYINPUT55), .A4(new_n579_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT109), .B1(new_n580_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n580_), .A2(new_n792_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n570_), .A2(new_n581_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n578_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n791_), .A2(new_n793_), .A3(new_n794_), .A4(new_n796_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT56), .B1(new_n797_), .B2(new_n589_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n786_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n477_), .B1(new_n473_), .B2(new_n469_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n469_), .B1(new_n471_), .B2(new_n465_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n468_), .A2(new_n802_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n474_), .A2(new_n477_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n593_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n657_), .B1(new_n800_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n785_), .B1(new_n806_), .B2(KEYINPUT57), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  INV_X1    g607(.A(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n797_), .A2(new_n589_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n809_), .B1(new_n814_), .B2(new_n786_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT110), .B(new_n808_), .C1(new_n815_), .C2(new_n657_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n806_), .A2(KEYINPUT57), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n804_), .A2(new_n592_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT111), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n804_), .A2(new_n820_), .A3(new_n592_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n799_), .B2(new_n798_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n814_), .A2(KEYINPUT58), .A3(new_n822_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n663_), .A3(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n807_), .A2(new_n816_), .A3(new_n817_), .A4(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n620_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n623_), .A2(new_n830_), .A3(new_n629_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT54), .B1(new_n622_), .B2(new_n478_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n784_), .B1(new_n829_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n559_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n836_), .A2(new_n826_), .B1(new_n806_), .B2(KEYINPUT57), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n808_), .B1(new_n815_), .B2(new_n657_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n621_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n831_), .A2(new_n832_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n783_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n844_), .B2(new_n783_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n835_), .A2(KEYINPUT59), .B1(new_n842_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n478_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G113gat), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n629_), .A2(G113gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n835_), .B2(new_n850_), .ZN(G1340gat));
  OAI21_X1  g650(.A(new_n846_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n597_), .B(new_n852_), .C1(new_n834_), .C2(new_n843_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G120gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n598_), .A2(KEYINPUT60), .ZN(new_n855_));
  MUX2_X1   g654(.A(new_n855_), .B(KEYINPUT60), .S(G120gat), .Z(new_n856_));
  NAND2_X1  g655(.A1(new_n834_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n854_), .A2(KEYINPUT113), .A3(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1341gat));
  AOI21_X1  g661(.A(G127gat), .B1(new_n834_), .B2(new_n621_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n621_), .A2(G127gat), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n864_), .B(KEYINPUT114), .Z(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n847_), .B2(new_n865_), .ZN(G1342gat));
  NAND2_X1  g665(.A1(new_n663_), .A2(G134gat), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT115), .Z(new_n868_));
  NAND2_X1  g667(.A1(new_n847_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n870_));
  AOI21_X1  g669(.A(G134gat), .B1(new_n834_), .B2(new_n657_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(new_n870_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n840_), .B1(new_n620_), .B2(new_n828_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT59), .B1(new_n874_), .B2(new_n784_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n875_), .A2(new_n852_), .A3(new_n868_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT116), .B1(new_n876_), .B2(new_n871_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n877_), .ZN(G1343gat));
  NAND3_X1  g677(.A1(new_n285_), .A2(new_n410_), .A3(new_n431_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n874_), .A2(new_n635_), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n478_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G141gat), .ZN(G1344gat));
  XNOR2_X1  g681(.A(KEYINPUT117), .B(G148gat), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n880_), .A2(new_n885_), .A3(new_n597_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n880_), .B2(new_n597_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n880_), .A2(new_n597_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT118), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n880_), .A2(new_n885_), .A3(new_n597_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n883_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n892_), .ZN(G1345gat));
  NAND2_X1  g692(.A1(new_n880_), .A2(new_n621_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(G162gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n880_), .A2(new_n897_), .A3(new_n657_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n880_), .A2(new_n663_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1347gat));
  NOR3_X1   g699(.A1(new_n442_), .A2(new_n285_), .A3(new_n431_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n410_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n478_), .B(new_n903_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G169gat), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n903_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n841_), .A2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n478_), .A3(new_n297_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n904_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n907_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n907_), .A2(new_n910_), .A3(KEYINPUT119), .A4(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1348gat));
  NAND2_X1  g715(.A1(new_n829_), .A2(new_n833_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n409_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n918_), .A2(new_n213_), .A3(new_n598_), .A4(new_n902_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G176gat), .B1(new_n909_), .B2(new_n597_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n920_), .A2(KEYINPUT120), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(KEYINPUT120), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n919_), .B1(new_n921_), .B2(new_n922_), .ZN(G1349gat));
  NAND2_X1  g722(.A1(new_n842_), .A2(new_n903_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n924_), .A2(new_n292_), .A3(new_n620_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n918_), .A2(new_n620_), .A3(new_n902_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n926_), .A2(KEYINPUT121), .ZN(new_n927_));
  AOI21_X1  g726(.A(G183gat), .B1(new_n926_), .B2(KEYINPUT121), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n925_), .B1(new_n927_), .B2(new_n928_), .ZN(G1350gat));
  NAND2_X1  g728(.A1(new_n657_), .A2(new_n293_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT122), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n909_), .A2(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n233_), .B1(new_n909_), .B2(new_n663_), .ZN(new_n933_));
  OR3_X1    g732(.A1(new_n932_), .A2(new_n933_), .A3(KEYINPUT123), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT123), .B1(new_n932_), .B2(new_n933_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1351gat));
  NAND3_X1  g735(.A1(new_n635_), .A2(new_n285_), .A3(new_n667_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n874_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n478_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g739(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT124), .B(G204gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n597_), .ZN(new_n943_));
  MUX2_X1   g742(.A(new_n941_), .B(new_n942_), .S(new_n943_), .Z(G1353gat));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n945_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n938_), .A2(new_n621_), .A3(new_n947_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n945_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n949_));
  XOR2_X1   g748(.A(new_n949_), .B(KEYINPUT126), .Z(new_n950_));
  XNOR2_X1  g749(.A(new_n948_), .B(new_n950_), .ZN(G1354gat));
  NAND2_X1  g750(.A1(new_n938_), .A2(new_n657_), .ZN(new_n952_));
  XOR2_X1   g751(.A(KEYINPUT127), .B(G218gat), .Z(new_n953_));
  NOR2_X1   g752(.A1(new_n559_), .A2(new_n953_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n952_), .A2(new_n953_), .B1(new_n938_), .B2(new_n954_), .ZN(G1355gat));
endmodule


