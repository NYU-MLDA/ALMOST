//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT85), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT24), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n216_), .B2(new_n212_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT77), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT23), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(KEYINPUT23), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n217_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT74), .ZN(new_n228_));
  INV_X1    g027(.A(G183gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT25), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(G183gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n228_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT75), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT76), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT26), .A4(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237_));
  INV_X1    g036(.A(G190gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(KEYINPUT76), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(KEYINPUT75), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT74), .B1(new_n231_), .B2(G183gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n233_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n223_), .A2(new_n218_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n229_), .B1(new_n238_), .B2(KEYINPUT75), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n234_), .A2(G190gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n247_));
  OAI221_X1 g046(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .C1(new_n247_), .C2(new_n223_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G169gat), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n227_), .A2(new_n243_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G197gat), .B(G204gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G211gat), .B(G218gat), .ZN(new_n254_));
  OAI211_X1 g053(.A(KEYINPUT21), .B(new_n253_), .C1(new_n254_), .C2(KEYINPUT81), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  INV_X1    g055(.A(G218gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G211gat), .ZN(new_n258_));
  INV_X1    g057(.A(G211gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G218gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT81), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n256_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(G197gat), .A2(G204gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G197gat), .A2(G204gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(new_n254_), .B2(KEYINPUT21), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n252_), .B(new_n255_), .C1(new_n263_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n259_), .A2(G218gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n257_), .A2(G211gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n256_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT81), .B1(new_n258_), .B2(new_n260_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n272_), .B(new_n266_), .C1(new_n273_), .C2(new_n256_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n252_), .B1(new_n274_), .B2(new_n255_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n251_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n211_), .B1(new_n276_), .B2(KEYINPUT20), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n255_), .B1(new_n263_), .B2(new_n267_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n223_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(new_n225_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT86), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT22), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(G169gat), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT22), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n286_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(KEYINPUT22), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(G169gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT86), .ZN(new_n294_));
  AOI21_X1  g093(.A(G176gat), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n215_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n295_), .A2(KEYINPUT87), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT87), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT86), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT86), .B1(new_n292_), .B2(new_n293_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n298_), .B1(new_n302_), .B2(new_n215_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n285_), .B1(new_n297_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n244_), .B1(new_n247_), .B2(new_n223_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n230_), .A2(new_n232_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT26), .B(G190gat), .ZN(new_n307_));
  AOI211_X1 g106(.A(new_n217_), .B(new_n305_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n279_), .B1(new_n304_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n277_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n276_), .A2(new_n211_), .A3(KEYINPUT20), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n210_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT87), .B1(new_n295_), .B2(new_n296_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n302_), .A2(new_n298_), .A3(new_n215_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n284_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n316_), .A2(new_n278_), .A3(new_n308_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n278_), .A2(KEYINPUT82), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n268_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT20), .B1(new_n319_), .B2(new_n251_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n317_), .A2(new_n320_), .A3(new_n209_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n207_), .B1(new_n313_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT88), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n278_), .B1(new_n316_), .B2(new_n308_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n319_), .B2(new_n251_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n324_), .B1(new_n326_), .B2(new_n211_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n312_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n209_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n321_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n206_), .A3(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n322_), .A2(new_n323_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT27), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n245_), .A2(new_n246_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n250_), .B1(new_n305_), .B2(new_n334_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n233_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n212_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(new_n214_), .C1(new_n281_), .C2(new_n225_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n335_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n268_), .B2(new_n318_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT85), .B1(new_n341_), .B2(new_n325_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n312_), .A3(new_n324_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n321_), .B1(new_n209_), .B2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(KEYINPUT88), .A3(new_n206_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n332_), .A2(new_n333_), .A3(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n342_), .A2(new_n210_), .A3(new_n312_), .A4(new_n324_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n269_), .A2(new_n275_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n325_), .B1(new_n349_), .B2(new_n340_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n304_), .A2(new_n279_), .A3(new_n309_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n210_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n347_), .B1(new_n348_), .B2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n311_), .A2(KEYINPUT94), .A3(new_n210_), .A4(new_n312_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n207_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(KEYINPUT27), .A3(new_n331_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n346_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G1gat), .B(G29gat), .Z(new_n359_));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G127gat), .B(G134gat), .Z(new_n365_));
  XOR2_X1   g164(.A(G113gat), .B(G120gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(KEYINPUT91), .B(KEYINPUT4), .Z(new_n369_));
  NAND2_X1  g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(KEYINPUT1), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n377_), .B2(KEYINPUT1), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n376_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT80), .B(new_n375_), .C1(new_n377_), .C2(KEYINPUT1), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n374_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n377_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n375_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n372_), .B(KEYINPUT3), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n370_), .B(KEYINPUT2), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n368_), .B(new_n369_), .C1(new_n382_), .C2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n389_), .B(KEYINPUT90), .Z(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n382_), .A2(new_n387_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT89), .B1(new_n392_), .B2(new_n367_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n368_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n368_), .B(KEYINPUT89), .C1(new_n382_), .C2(new_n387_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n391_), .B1(new_n397_), .B2(KEYINPUT4), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n390_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n364_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n401_), .B(new_n363_), .C1(new_n403_), .C2(new_n391_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT29), .B1(new_n382_), .B2(new_n387_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n278_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(G228gat), .A3(G233gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G228gat), .A2(G233gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n349_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n408_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n392_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT28), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT28), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n392_), .A2(new_n419_), .A3(new_n416_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G22gat), .B(G50gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n420_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n421_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n411_), .A2(new_n413_), .A3(new_n408_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n415_), .A2(new_n422_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n415_), .A2(new_n428_), .A3(new_n426_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n414_), .A2(KEYINPUT83), .B1(new_n425_), .B2(new_n422_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n406_), .A2(new_n427_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n427_), .A2(new_n406_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n434_), .B(KEYINPUT78), .Z(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT30), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n251_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT31), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT79), .B1(new_n367_), .B2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n440_), .B2(new_n367_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G15gat), .B(G43gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n439_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NOR4_X1   g245(.A1(new_n358_), .A2(new_n405_), .A3(new_n433_), .A4(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n400_), .A2(new_n404_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n355_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n448_), .B1(KEYINPUT95), .B2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n329_), .A2(new_n330_), .A3(new_n449_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n344_), .A2(KEYINPUT93), .A3(new_n449_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n449_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n455_), .A2(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n332_), .A2(new_n345_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n390_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n388_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n403_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n463_), .A2(new_n363_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n404_), .A2(KEYINPUT33), .ZN(new_n466_));
  INV_X1    g265(.A(new_n398_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT33), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n401_), .A4(new_n363_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n465_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n452_), .A2(new_n459_), .B1(new_n460_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n405_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OAI22_X1  g272(.A1(new_n471_), .A2(new_n433_), .B1(new_n473_), .B2(new_n358_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n447_), .B1(new_n474_), .B2(new_n446_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT65), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT9), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT64), .B(G92gat), .ZN(new_n478_));
  INV_X1    g277(.A(G85gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G92gat), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n477_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n476_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n481_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n482_), .B1(KEYINPUT65), .B2(new_n485_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT10), .B(G99gat), .Z(new_n492_));
  AOI21_X1  g291(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G85gat), .B(G92gat), .Z(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  INV_X1    g294(.A(G99gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n491_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n494_), .B1(new_n490_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT8), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n500_), .A2(KEYINPUT8), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n487_), .A2(new_n493_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G29gat), .B(G36gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT35), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT34), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n503_), .A2(new_n506_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n507_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n493_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT66), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n502_), .A2(new_n501_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT66), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n517_), .B(new_n493_), .C1(new_n484_), .C2(new_n486_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n506_), .B(KEYINPUT15), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n511_), .A2(new_n513_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n513_), .B1(new_n511_), .B2(new_n521_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G190gat), .B(G218gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G134gat), .B(G162gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT36), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  NOR4_X1   g330(.A1(new_n523_), .A2(new_n524_), .A3(KEYINPUT36), .A4(new_n528_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n537_));
  XOR2_X1   g336(.A(G71gat), .B(G78gat), .Z(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n537_), .A2(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n516_), .B2(new_n514_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n534_), .B1(new_n542_), .B2(KEYINPUT12), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n544_));
  OAI211_X1 g343(.A(KEYINPUT67), .B(new_n544_), .C1(new_n503_), .C2(new_n541_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT68), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G230gat), .A2(G233gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n539_), .A2(KEYINPUT12), .A3(new_n540_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n519_), .A2(new_n550_), .B1(new_n503_), .B2(new_n541_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .A4(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n548_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n503_), .A2(new_n541_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(new_n542_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n551_), .A2(new_n543_), .A3(new_n545_), .A4(new_n548_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT68), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G120gat), .B(G148gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT70), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n558_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n552_), .A2(new_n555_), .A3(new_n557_), .A4(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT13), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n570_), .A3(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573_));
  INV_X1    g372(.A(G8gat), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G1gat), .B(G8gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n541_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583_));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n582_), .A2(new_n583_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(KEYINPUT17), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n582_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n578_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n520_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT72), .Z(new_n595_));
  NAND2_X1  g394(.A1(G229gat), .A2(G233gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n506_), .B(KEYINPUT71), .Z(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n578_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n578_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n595_), .A2(new_n599_), .B1(new_n600_), .B2(new_n597_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT73), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G169gat), .B(G197gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n605_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n572_), .A2(new_n592_), .A3(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n475_), .A2(new_n533_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n202_), .B1(new_n610_), .B2(new_n405_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT97), .Z(new_n612_));
  INV_X1    g411(.A(new_n608_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n572_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n533_), .B(KEYINPUT37), .Z(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n592_), .ZN(new_n616_));
  NOR4_X1   g415(.A1(new_n475_), .A2(new_n613_), .A3(new_n614_), .A4(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  AOI21_X1  g417(.A(G1gat), .B1(new_n618_), .B2(KEYINPUT96), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n405_), .A3(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n618_), .A2(KEYINPUT96), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n612_), .A2(new_n622_), .ZN(G1324gat));
  AOI21_X1  g422(.A(new_n574_), .B1(new_n610_), .B2(new_n358_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT39), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n617_), .A2(new_n574_), .A3(new_n358_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g427(.A(G15gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n610_), .B2(new_n445_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n617_), .A2(new_n629_), .A3(new_n445_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n610_), .B2(new_n433_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT42), .Z(new_n636_));
  NAND3_X1  g435(.A1(new_n617_), .A2(new_n634_), .A3(new_n433_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1327gat));
  OAI21_X1  g437(.A(KEYINPUT43), .B1(new_n475_), .B2(new_n615_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n451_), .A2(KEYINPUT95), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n457_), .A2(new_n458_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n455_), .A2(new_n456_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n640_), .A2(new_n405_), .A3(new_n641_), .A4(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n323_), .B1(new_n344_), .B2(new_n206_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n331_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n345_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n470_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n433_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n472_), .A2(new_n346_), .A3(new_n357_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n446_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n358_), .A2(new_n433_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n446_), .A2(new_n405_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n533_), .B(KEYINPUT37), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n639_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n571_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n570_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n591_), .B(new_n608_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT44), .B1(new_n659_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n667_), .B(new_n664_), .C1(new_n639_), .C2(new_n658_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n448_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n533_), .A2(new_n591_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n614_), .A2(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n655_), .A2(new_n608_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n675_), .A2(G29gat), .A3(new_n448_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n676_), .ZN(G1328gat));
  NAND2_X1  g476(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n678_));
  NOR2_X1   g477(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n679_));
  AOI21_X1  g478(.A(G36gat), .B1(new_n346_), .B2(new_n357_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n655_), .A2(new_n608_), .A3(new_n673_), .A4(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT100), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT100), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT45), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n682_), .A2(new_n686_), .A3(new_n683_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n679_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT99), .B1(new_n669_), .B2(new_n358_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n656_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT43), .B(new_n615_), .C1(new_n651_), .C2(new_n654_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n665_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n667_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n665_), .B(KEYINPUT44), .C1(new_n690_), .C2(new_n691_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n693_), .A2(KEYINPUT99), .A3(new_n358_), .A4(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G36gat), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n678_), .B(new_n688_), .C1(new_n689_), .C2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n693_), .A2(new_n358_), .A3(new_n694_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(G36gat), .A3(new_n695_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n678_), .B1(new_n702_), .B2(new_n688_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n698_), .A2(new_n703_), .ZN(G1329gat));
  NAND3_X1  g503(.A1(new_n669_), .A2(G43gat), .A3(new_n445_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n675_), .A2(new_n446_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(G43gat), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g507(.A(new_n433_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G50gat), .B1(new_n670_), .B2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(G50gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT102), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n675_), .B2(new_n712_), .ZN(G1331gat));
  NOR2_X1   g512(.A1(new_n616_), .A2(new_n572_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT103), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n655_), .A2(new_n613_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n405_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n533_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n572_), .A2(new_n591_), .A3(new_n608_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n655_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT104), .Z(new_n722_));
  NOR2_X1   g521(.A1(new_n448_), .A2(KEYINPUT105), .ZN(new_n723_));
  MUX2_X1   g522(.A(KEYINPUT105), .B(new_n723_), .S(G57gat), .Z(new_n724_));
  AOI21_X1  g523(.A(new_n718_), .B1(new_n722_), .B2(new_n724_), .ZN(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n717_), .A2(new_n726_), .A3(new_n358_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n722_), .A2(new_n358_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G64gat), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n717_), .A2(new_n733_), .A3(new_n445_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n722_), .A2(new_n445_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G71gat), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(KEYINPUT49), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(KEYINPUT49), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1334gat));
  INV_X1    g538(.A(G78gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n717_), .A2(new_n740_), .A3(new_n433_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n722_), .A2(new_n433_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G78gat), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT50), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT50), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1335gat));
  NOR3_X1   g545(.A1(new_n716_), .A2(new_n572_), .A3(new_n672_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n479_), .A3(new_n405_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n572_), .A2(new_n592_), .A3(new_n608_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n659_), .A2(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n405_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n751_), .B2(new_n479_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT106), .ZN(G1336gat));
  AOI21_X1  g552(.A(G92gat), .B1(new_n747_), .B2(new_n358_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n478_), .B1(new_n346_), .B2(new_n357_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT107), .Z(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n750_), .B2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT108), .Z(G1337gat));
  NAND3_X1  g557(.A1(new_n747_), .A2(new_n445_), .A3(new_n492_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n750_), .A2(new_n445_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n496_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n659_), .A2(new_n433_), .A3(new_n749_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(G106gat), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n763_), .A3(G106gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n709_), .A2(G106gat), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n765_), .A2(new_n766_), .B1(new_n747_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n769_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1339gat));
  XOR2_X1   g574(.A(KEYINPUT114), .B(G113gat), .Z(new_n776_));
  NAND2_X1  g575(.A1(new_n608_), .A2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT115), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n615_), .A2(new_n572_), .A3(new_n592_), .A4(new_n613_), .ZN(new_n779_));
  XOR2_X1   g578(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n779_), .B(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n608_), .A2(new_n567_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n551_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n553_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(new_n556_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n552_), .A2(new_n786_), .A3(new_n557_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n565_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n792_), .B(new_n564_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n783_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n596_), .B1(new_n598_), .B2(new_n578_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n595_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n605_), .B1(new_n600_), .B2(new_n596_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n601_), .A2(new_n605_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n568_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n794_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n719_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n798_), .A2(new_n567_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT112), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n798_), .A2(new_n567_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n615_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n552_), .A2(new_n786_), .A3(new_n557_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n565_), .B1(new_n812_), .B2(new_n787_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n792_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n565_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n814_), .A2(new_n815_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n811_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n533_), .B1(new_n794_), .B2(new_n799_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n803_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n782_), .B1(new_n821_), .B2(new_n591_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n652_), .A2(new_n405_), .A3(new_n445_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n657_), .B1(new_n816_), .B2(KEYINPUT58), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n809_), .A2(new_n810_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n826_), .A2(new_n827_), .B1(new_n819_), .B2(KEYINPUT57), .ZN(new_n828_));
  INV_X1    g627(.A(new_n820_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n591_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n782_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n824_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT59), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n778_), .B1(new_n825_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(new_n608_), .A3(new_n833_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n835_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n835_), .B(KEYINPUT116), .C1(new_n839_), .C2(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1340gat));
  NAND2_X1  g644(.A1(new_n832_), .A2(new_n833_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n572_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n847_), .B(new_n849_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n823_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n832_), .A2(KEYINPUT59), .A3(new_n833_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n572_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854_));
  OAI21_X1  g653(.A(G120gat), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n825_), .A2(new_n834_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n856_), .A2(KEYINPUT117), .A3(new_n572_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n850_), .B1(new_n855_), .B2(new_n857_), .ZN(G1341gat));
  OAI21_X1  g657(.A(G127gat), .B1(new_n856_), .B2(new_n591_), .ZN(new_n859_));
  OR3_X1    g658(.A1(new_n846_), .A2(G127gat), .A3(new_n591_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1342gat));
  XOR2_X1   g660(.A(KEYINPUT118), .B(G134gat), .Z(new_n862_));
  NOR3_X1   g661(.A1(new_n856_), .A2(new_n615_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(G134gat), .B1(new_n847_), .B2(new_n533_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1343gat));
  NOR4_X1   g664(.A1(new_n358_), .A2(new_n709_), .A3(new_n448_), .A4(new_n445_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n832_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n608_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n614_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n867_), .A2(new_n591_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT61), .B(G155gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  INV_X1    g674(.A(G162gat), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n867_), .A2(new_n876_), .A3(new_n615_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n867_), .B2(new_n719_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n878_), .A2(KEYINPUT119), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(KEYINPUT119), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n877_), .B1(new_n879_), .B2(new_n880_), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n358_), .A2(new_n653_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT120), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n822_), .A2(new_n433_), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n608_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G169gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n887_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n885_), .A2(G169gat), .A3(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n300_), .A2(new_n301_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n888_), .B(new_n890_), .C1(new_n891_), .C2(new_n885_), .ZN(G1348gat));
  NAND2_X1  g691(.A1(new_n884_), .A2(new_n614_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g693(.A1(new_n884_), .A2(new_n592_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(G183gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n306_), .B1(KEYINPUT122), .B2(G183gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n895_), .B2(new_n898_), .ZN(G1350gat));
  INV_X1    g698(.A(new_n884_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G190gat), .B1(new_n900_), .B2(new_n615_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n884_), .A2(new_n307_), .A3(new_n533_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1351gat));
  NAND3_X1  g702(.A1(new_n472_), .A2(KEYINPUT123), .A3(new_n446_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n358_), .ZN(new_n905_));
  AOI21_X1  g704(.A(KEYINPUT123), .B1(new_n472_), .B2(new_n446_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n832_), .A2(new_n608_), .A3(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n908_), .A2(new_n909_), .A3(KEYINPUT125), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT125), .B1(new_n908_), .B2(new_n909_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n909_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G197gat), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n910_), .A2(G197gat), .A3(new_n911_), .A4(new_n913_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1352gat));
  NOR3_X1   g716(.A1(new_n822_), .A2(new_n906_), .A3(new_n905_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n614_), .ZN(new_n919_));
  INV_X1    g718(.A(G204gat), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(KEYINPUT126), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n919_), .B(new_n921_), .ZN(G1353gat));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n591_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n918_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n923_), .B1(new_n918_), .B2(new_n924_), .ZN(new_n927_));
  OAI22_X1  g726(.A1(new_n926_), .A2(new_n927_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  INV_X1    g727(.A(new_n927_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(new_n930_), .A3(new_n925_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n928_), .A2(new_n931_), .ZN(G1354gat));
  NAND3_X1  g731(.A1(new_n918_), .A2(new_n257_), .A3(new_n533_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n918_), .A2(new_n657_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(new_n257_), .ZN(G1355gat));
endmodule


