//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT36), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G85gat), .A3(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G85gat), .B(G92gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n206_), .B2(new_n204_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT65), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  AND2_X1   g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT10), .B(G99gat), .Z(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n208_), .A2(new_n216_), .A3(new_n217_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n213_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n209_), .A2(KEYINPUT65), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(KEYINPUT66), .A3(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT7), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n224_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n206_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n222_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  AOI211_X1 g034(.A(KEYINPUT8), .B(new_n206_), .C1(new_n216_), .C2(new_n232_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n221_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G29gat), .B(G36gat), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n238_), .A2(KEYINPUT70), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(KEYINPUT70), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G43gat), .B(G50gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n239_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n245_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n246_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n237_), .A2(new_n247_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G232gat), .A2(G233gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT34), .Z(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n254_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n221_), .B(new_n248_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n251_), .A2(new_n256_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G190gat), .B(G218gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G134gat), .B(G162gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT73), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(KEYINPUT72), .A3(new_n257_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n251_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT72), .B1(new_n258_), .B2(new_n257_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n263_), .B(new_n255_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n258_), .A2(new_n257_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(new_n264_), .A3(new_n251_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n263_), .B1(new_n272_), .B2(new_n255_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n259_), .B(new_n262_), .C1(new_n268_), .C2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(KEYINPUT74), .B(new_n259_), .C1(new_n268_), .C2(new_n273_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n262_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n203_), .A2(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n275_), .A2(new_n203_), .A3(new_n276_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n202_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT37), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(new_n203_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n275_), .A2(new_n203_), .A3(new_n276_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(new_n202_), .A3(KEYINPUT37), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G15gat), .B(G22gat), .ZN(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n290_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n293_), .A2(new_n294_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G8gat), .ZN(new_n297_));
  OR3_X1    g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n297_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G231gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G57gat), .B(G64gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT11), .ZN(new_n304_));
  XOR2_X1   g103(.A(G71gat), .B(G78gat), .Z(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n303_), .A2(KEYINPUT11), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n304_), .A2(new_n305_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n302_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(new_n311_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT77), .ZN(new_n315_));
  XOR2_X1   g114(.A(G127gat), .B(G155gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G183gat), .B(G211gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(KEYINPUT77), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n315_), .A2(KEYINPUT17), .A3(new_n321_), .A4(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n314_), .A2(KEYINPUT79), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n314_), .A2(KEYINPUT79), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n320_), .B(KEYINPUT17), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n289_), .A2(KEYINPUT80), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n237_), .A2(new_n311_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n221_), .B(new_n310_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n334_), .B(new_n336_), .C1(new_n332_), .C2(new_n331_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n335_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT68), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT68), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n333_), .A2(new_n340_), .A3(new_n335_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n237_), .B2(new_n311_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n237_), .A2(new_n342_), .A3(new_n311_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n339_), .B(new_n341_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n337_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G120gat), .B(G148gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT5), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G176gat), .B(G204gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT13), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(KEYINPUT13), .A3(new_n352_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n288_), .B2(new_n328_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n330_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT81), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n300_), .B(new_n248_), .Z(new_n362_));
  NAND2_X1  g161(.A1(G229gat), .A2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n250_), .A2(new_n300_), .A3(new_n247_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n248_), .A2(new_n299_), .A3(new_n298_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G113gat), .B(G141gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G169gat), .B(G197gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n369_), .A2(new_n370_), .A3(new_n374_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n376_), .A2(KEYINPUT83), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT83), .B1(new_n376_), .B2(new_n377_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G155gat), .B(G162gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT92), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n381_), .A2(KEYINPUT92), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G141gat), .A2(G148gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT2), .ZN(new_n385_));
  INV_X1    g184(.A(G141gat), .ZN(new_n386_));
  INV_X1    g185(.A(G148gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT91), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n388_), .A2(new_n389_), .A3(KEYINPUT3), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n382_), .B(new_n383_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n388_), .A2(new_n384_), .A3(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(KEYINPUT1), .B2(new_n381_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT93), .ZN(new_n398_));
  XOR2_X1   g197(.A(G127gat), .B(G134gat), .Z(new_n399_));
  XNOR2_X1  g198(.A(G113gat), .B(G120gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n397_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n401_), .A2(KEYINPUT101), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(KEYINPUT101), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  MUX2_X1   g209(.A(new_n402_), .B(new_n407_), .S(KEYINPUT4), .Z(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(new_n409_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G85gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT0), .B(G57gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n414_), .B(new_n415_), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n412_), .A2(new_n416_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT103), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n419_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT103), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n417_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G197gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G204gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT96), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n425_), .A2(G204gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT95), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(KEYINPUT95), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT21), .ZN(new_n433_));
  XOR2_X1   g232(.A(G211gat), .B(G218gat), .Z(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(KEYINPUT97), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n432_), .B(new_n435_), .C1(KEYINPUT97), .C2(new_n434_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n429_), .A2(new_n426_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(KEYINPUT21), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n432_), .B2(KEYINPUT21), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(KEYINPUT89), .B(G176gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT22), .B(G169gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G169gat), .A2(G176gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n444_), .B(KEYINPUT87), .Z(new_n445_));
  AND2_X1   g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G183gat), .A2(G190gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT23), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(G183gat), .B2(G190gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n444_), .A2(KEYINPUT24), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT100), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G169gat), .A2(G176gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT86), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT26), .B(G190gat), .ZN(new_n456_));
  INV_X1    g255(.A(G183gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT25), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n457_), .A2(KEYINPUT25), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n453_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n460_), .B(new_n448_), .C1(KEYINPUT24), .C2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n450_), .B1(new_n455_), .B2(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n440_), .A2(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n464_), .A2(KEYINPUT20), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G226gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT85), .B(G190gat), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n469_), .A2(new_n457_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n448_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n446_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n448_), .B1(new_n454_), .B2(KEYINPUT24), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n458_), .B(KEYINPUT84), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT26), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n476_), .B(new_n459_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n445_), .A2(KEYINPUT24), .A3(new_n454_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n475_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n473_), .A2(new_n474_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n472_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n440_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n465_), .A2(new_n468_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G8gat), .B(G36gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT18), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G64gat), .B(G92gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n440_), .A2(new_n463_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(KEYINPUT20), .C1(new_n484_), .C2(new_n440_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n468_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n486_), .A2(new_n490_), .A3(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n492_), .A2(new_n493_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n465_), .A2(KEYINPUT102), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n464_), .A2(KEYINPUT20), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT102), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n485_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n496_), .B1(new_n501_), .B2(new_n493_), .ZN(new_n502_));
  OAI211_X1 g301(.A(KEYINPUT27), .B(new_n495_), .C1(new_n502_), .C2(new_n490_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n486_), .A2(new_n494_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n490_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n495_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT27), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G228gat), .A2(G233gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n397_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT29), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n512_), .B(new_n440_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n440_), .B1(new_n403_), .B2(new_n515_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G228gat), .A3(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G78gat), .B(G106gat), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT98), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G22gat), .B(G50gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n398_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT28), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n525_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT28), .B1(new_n398_), .B2(KEYINPUT29), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n514_), .A2(new_n527_), .A3(new_n515_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n524_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n529_), .A2(KEYINPUT94), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT94), .B1(new_n529_), .B2(new_n532_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n522_), .B(new_n523_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n532_), .B(new_n529_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G227gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(G71gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(G99gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n484_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(new_n401_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G15gat), .B(G43gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT90), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT30), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT31), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n543_), .B(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n522_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT98), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n537_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n548_), .B1(new_n537_), .B2(new_n550_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n424_), .B(new_n511_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n537_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n550_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n490_), .A2(KEYINPUT32), .ZN(new_n557_));
  MUX2_X1   g356(.A(new_n502_), .B(new_n504_), .S(new_n557_), .Z(new_n558_));
  OAI21_X1  g357(.A(new_n558_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n416_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n411_), .B2(new_n408_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n507_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT33), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n412_), .A2(new_n564_), .A3(new_n416_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n563_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n559_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n548_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n556_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n380_), .B1(new_n553_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT81), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n330_), .A2(new_n572_), .A3(new_n357_), .A4(new_n359_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n424_), .A2(G1gat), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n361_), .A2(new_n571_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT104), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT104), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(KEYINPUT38), .A3(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n376_), .A2(new_n377_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n357_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT105), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n329_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n286_), .B1(new_n553_), .B2(new_n570_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n583_), .A2(KEYINPUT106), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(KEYINPUT106), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n582_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(G1gat), .B1(new_n587_), .B2(new_n424_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n578_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT38), .B1(new_n576_), .B2(new_n577_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(G1324gat));
  AOI211_X1 g390(.A(new_n511_), .B(new_n582_), .C1(new_n585_), .C2(new_n584_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT39), .B1(new_n592_), .B2(new_n292_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n594_), .B(G8gat), .C1(new_n587_), .C2(new_n511_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n361_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n292_), .A3(new_n510_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT40), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n596_), .A2(KEYINPUT40), .A3(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1325gat));
  INV_X1    g402(.A(G15gat), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n586_), .B2(new_n548_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT41), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n597_), .A2(new_n604_), .A3(new_n548_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1326gat));
  INV_X1    g407(.A(G22gat), .ZN(new_n609_));
  INV_X1    g408(.A(new_n556_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n586_), .B2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT42), .Z(new_n612_));
  NAND3_X1  g411(.A1(new_n597_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(G1327gat));
  NAND2_X1  g413(.A1(new_n553_), .A2(new_n570_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n288_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(KEYINPUT43), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(KEYINPUT43), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n328_), .B(new_n581_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n424_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n616_), .B(KEYINPUT43), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n623_), .A2(KEYINPUT44), .A3(new_n328_), .A4(new_n581_), .ZN(new_n624_));
  AND4_X1   g423(.A1(G29gat), .A2(new_n621_), .A3(new_n622_), .A4(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n286_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n329_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n571_), .A2(new_n357_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n622_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n625_), .A2(new_n629_), .ZN(G1328gat));
  NAND3_X1  g429(.A1(new_n621_), .A2(new_n510_), .A3(new_n624_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G36gat), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n511_), .A2(KEYINPUT107), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n511_), .A2(KEYINPUT107), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(G36gat), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n628_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT45), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n632_), .B(new_n638_), .C1(KEYINPUT108), .C2(KEYINPUT46), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1329gat));
  NAND4_X1  g442(.A1(new_n621_), .A2(new_n624_), .A3(G43gat), .A4(new_n548_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT109), .B(G43gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n628_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(new_n569_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(G1330gat));
  AND4_X1   g449(.A1(G50gat), .A2(new_n621_), .A3(new_n610_), .A4(new_n624_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G50gat), .B1(new_n628_), .B2(new_n610_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1331gat));
  NAND2_X1  g452(.A1(new_n584_), .A2(new_n585_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n380_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n357_), .A2(new_n328_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G57gat), .B1(new_n657_), .B2(new_n424_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n330_), .A2(new_n359_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n357_), .A2(new_n579_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n615_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n424_), .A2(G57gat), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n658_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT111), .Z(G1332gat));
  OAI21_X1  g465(.A(G64gat), .B1(new_n657_), .B2(new_n635_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT48), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT48), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n635_), .A2(G64gat), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT112), .Z(new_n671_));
  OAI22_X1  g470(.A1(new_n668_), .A2(new_n669_), .B1(new_n662_), .B2(new_n671_), .ZN(G1333gat));
  INV_X1    g471(.A(new_n662_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n539_), .A3(new_n548_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G71gat), .B1(new_n657_), .B2(new_n569_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT49), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT49), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n674_), .B1(new_n676_), .B2(new_n677_), .ZN(G1334gat));
  INV_X1    g477(.A(G78gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n673_), .A2(new_n679_), .A3(new_n610_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n657_), .A2(new_n556_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n679_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n683_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n684_), .B2(new_n685_), .ZN(G1335gat));
  OAI211_X1 g485(.A(new_n328_), .B(new_n660_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G85gat), .B1(new_n687_), .B2(new_n424_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n661_), .A2(new_n627_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n424_), .A2(G85gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(G1336gat));
  INV_X1    g490(.A(G92gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n692_), .B1(new_n689_), .B2(new_n511_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT114), .Z(new_n694_));
  NOR3_X1   g493(.A1(new_n687_), .A2(new_n692_), .A3(new_n635_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1337gat));
  OAI21_X1  g495(.A(G99gat), .B1(new_n687_), .B2(new_n569_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n689_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n218_), .A3(new_n548_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g500(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n702_));
  OAI21_X1  g501(.A(G106gat), .B1(new_n687_), .B2(new_n556_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(G106gat), .B(new_n704_), .C1(new_n687_), .C2(new_n556_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n689_), .A2(G106gat), .A3(new_n556_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n702_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n702_), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n709_), .B(new_n712_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1339gat));
  AND4_X1   g513(.A1(new_n356_), .A2(new_n355_), .A3(new_n329_), .A4(new_n380_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n281_), .A2(new_n287_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT54), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT54), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n281_), .A2(new_n287_), .A3(new_n718_), .A4(new_n715_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n362_), .A2(new_n363_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n366_), .A2(new_n367_), .A3(new_n364_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n375_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n369_), .A2(new_n374_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n353_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n579_), .A2(new_n351_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT55), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n333_), .B1(new_n344_), .B2(new_n343_), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n345_), .A2(new_n728_), .B1(new_n336_), .B2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT117), .B1(new_n345_), .B2(new_n728_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n333_), .A2(new_n340_), .A3(new_n335_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n343_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n237_), .A2(new_n342_), .A3(new_n311_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT117), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(KEYINPUT55), .A4(new_n339_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n730_), .A2(new_n731_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n350_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT56), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n727_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT118), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n726_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n727_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n738_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT56), .B1(new_n738_), .B2(new_n350_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n746_), .B(new_n744_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n626_), .B1(new_n745_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n726_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(KEYINPUT118), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n286_), .B1(new_n756_), .B2(new_n749_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT57), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n741_), .A2(new_n742_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n351_), .A2(new_n725_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n759_), .A2(new_n760_), .A3(KEYINPUT58), .A4(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT58), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT58), .B(new_n761_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT120), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n288_), .A2(new_n762_), .A3(new_n765_), .A4(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n753_), .A2(new_n758_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n720_), .B1(new_n769_), .B2(new_n328_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n424_), .A2(new_n510_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n551_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(KEYINPUT59), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT122), .B1(new_n770_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT122), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n767_), .A2(new_n762_), .A3(new_n765_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n288_), .A2(new_n777_), .B1(new_n757_), .B2(KEYINPUT57), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n329_), .B1(new_n778_), .B2(new_n753_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n776_), .B(new_n773_), .C1(new_n779_), .C2(new_n720_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n775_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n751_), .A2(KEYINPUT119), .A3(new_n752_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n757_), .B2(KEYINPUT57), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n778_), .A2(new_n782_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n720_), .B1(new_n785_), .B2(new_n328_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT59), .B1(new_n786_), .B2(new_n772_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n781_), .A2(new_n655_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n790_));
  OR3_X1    g589(.A1(new_n786_), .A2(new_n790_), .A3(new_n772_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n786_), .B2(new_n772_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n579_), .A2(new_n789_), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n788_), .A2(new_n789_), .B1(new_n793_), .B2(new_n794_), .ZN(G1340gat));
  INV_X1    g594(.A(new_n357_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n781_), .A2(new_n796_), .A3(new_n787_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT123), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n781_), .A2(new_n787_), .A3(KEYINPUT123), .A4(new_n796_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(G120gat), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT60), .ZN(new_n802_));
  AOI21_X1  g601(.A(G120gat), .B1(new_n796_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n802_), .B2(G120gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n791_), .A2(new_n792_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n805_), .ZN(G1341gat));
  NAND3_X1  g605(.A1(new_n781_), .A2(new_n329_), .A3(new_n787_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G127gat), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n328_), .A2(G127gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n793_), .B2(new_n809_), .ZN(G1342gat));
  NAND3_X1  g609(.A1(new_n781_), .A2(new_n288_), .A3(new_n787_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G134gat), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n626_), .A2(G134gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n793_), .B2(new_n813_), .ZN(G1343gat));
  INV_X1    g613(.A(new_n552_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n786_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n635_), .A2(new_n622_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n579_), .A3(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n796_), .A3(new_n818_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g621(.A1(new_n816_), .A2(new_n329_), .A3(new_n818_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT61), .B(G155gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1346gat));
  INV_X1    g624(.A(G162gat), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n816_), .A2(new_n826_), .A3(new_n286_), .A4(new_n818_), .ZN(new_n827_));
  NOR4_X1   g626(.A1(new_n786_), .A2(new_n289_), .A3(new_n815_), .A4(new_n817_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n827_), .B(KEYINPUT124), .C1(new_n826_), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1347gat));
  NOR2_X1   g632(.A1(new_n635_), .A2(new_n622_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n548_), .A3(new_n579_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT125), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n770_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n556_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(G169gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT62), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n834_), .A2(new_n551_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n838_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n442_), .A3(new_n579_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n845_), .ZN(G1348gat));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n796_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n786_), .A2(new_n610_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n834_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n569_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n850_), .A2(G176gat), .A3(new_n796_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n847_), .A2(new_n441_), .B1(new_n848_), .B2(new_n851_), .ZN(G1349gat));
  NAND3_X1  g651(.A1(new_n848_), .A2(new_n329_), .A3(new_n850_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n328_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n853_), .A2(new_n457_), .B1(new_n844_), .B2(new_n854_), .ZN(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n843_), .B2(new_n289_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n286_), .A2(new_n456_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n843_), .B2(new_n857_), .ZN(G1351gat));
  NAND3_X1  g657(.A1(new_n816_), .A2(new_n579_), .A3(new_n834_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT126), .B(G197gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n859_), .B(new_n860_), .Z(G1352gat));
  NAND3_X1  g660(.A1(new_n816_), .A2(new_n796_), .A3(new_n834_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g662(.A1(new_n816_), .A2(new_n329_), .A3(new_n834_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  AND2_X1   g664(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n864_), .B2(new_n865_), .ZN(G1354gat));
  INV_X1    g667(.A(G218gat), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n816_), .A2(new_n869_), .A3(new_n286_), .A4(new_n834_), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n786_), .A2(new_n289_), .A3(new_n815_), .A4(new_n849_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT127), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n870_), .B(KEYINPUT127), .C1(new_n869_), .C2(new_n871_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1355gat));
endmodule


