//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  INV_X1    g006(.A(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT9), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G85gat), .A3(G92gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n202_), .B1(new_n212_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n219_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n221_), .A2(KEYINPUT65), .A3(new_n206_), .A4(new_n211_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT7), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n214_), .A2(KEYINPUT66), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT6), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n213_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n227_), .A2(new_n229_), .A3(new_n213_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n226_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n209_), .A2(new_n210_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n224_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n215_), .A2(new_n218_), .ZN(new_n238_));
  AOI211_X1 g037(.A(KEYINPUT8), .B(new_n235_), .C1(new_n226_), .C2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n223_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT73), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G43gat), .B(G50gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n242_), .A2(KEYINPUT73), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(KEYINPUT73), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n244_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n246_), .A2(KEYINPUT15), .A3(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(new_n241_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT34), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(KEYINPUT35), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(KEYINPUT35), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT75), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n256_), .A2(KEYINPUT75), .A3(new_n261_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n251_), .B(new_n259_), .C1(new_n255_), .C2(new_n241_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G190gat), .B(G218gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G134gat), .B(G162gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(KEYINPUT36), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT76), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT37), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n264_), .A2(new_n275_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n270_), .A2(KEYINPUT36), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n276_), .A2(new_n278_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n271_), .B(new_n274_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n272_), .A2(new_n273_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n276_), .B(new_n278_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n282_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n284_), .A2(new_n271_), .A3(new_n274_), .A4(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT14), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT77), .B(G8gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n289_), .B2(G1gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT78), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G15gat), .B(G22gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G8gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G57gat), .B(G64gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n300_));
  XOR2_X1   g099(.A(G71gat), .B(G78gat), .Z(new_n301_));
  OR2_X1    g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n301_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G231gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n298_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G127gat), .B(G155gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT16), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G183gat), .B(G211gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT17), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT79), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n308_), .B(KEYINPUT80), .Z(new_n316_));
  OR2_X1    g115(.A1(new_n312_), .A2(KEYINPUT17), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n313_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n318_), .A2(KEYINPUT81), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(KEYINPUT81), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n315_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n287_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT69), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n226_), .A2(new_n238_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(new_n224_), .A3(new_n236_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n227_), .A2(new_n229_), .A3(new_n213_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n213_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n235_), .B1(new_n328_), .B2(new_n226_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n325_), .B1(new_n329_), .B2(new_n224_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n305_), .B1(new_n330_), .B2(new_n223_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n323_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n305_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n240_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n332_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(KEYINPUT69), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n331_), .A2(KEYINPUT12), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n305_), .B(new_n223_), .C1(new_n237_), .C2(new_n239_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G230gat), .A2(G233gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT64), .Z(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n333_), .A2(new_n337_), .A3(new_n338_), .A4(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT70), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n332_), .B1(new_n240_), .B2(new_n334_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n346_), .A2(KEYINPUT69), .B1(new_n331_), .B2(KEYINPUT12), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n347_), .A2(KEYINPUT70), .A3(new_n333_), .A4(new_n342_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n341_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n339_), .A2(KEYINPUT67), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n335_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n339_), .A2(KEYINPUT67), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n349_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n345_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G120gat), .B(G148gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT5), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G176gat), .B(G204gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT71), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n358_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n345_), .A2(new_n348_), .A3(new_n353_), .A4(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n365_));
  OR2_X1    g164(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n364_), .A2(new_n366_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G155gat), .B(G162gat), .Z(new_n371_));
  INV_X1    g170(.A(KEYINPUT1), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374_));
  INV_X1    g173(.A(G141gat), .ZN(new_n375_));
  INV_X1    g174(.A(G148gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n373_), .A2(new_n374_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT88), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n374_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n381_), .B(new_n382_), .C1(new_n384_), .C2(KEYINPUT2), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n384_), .A2(KEYINPUT2), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n371_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n379_), .A2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G127gat), .B(G134gat), .Z(new_n389_));
  XOR2_X1   g188(.A(G113gat), .B(G120gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n379_), .A2(new_n387_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n392_), .A2(KEYINPUT4), .A3(new_n395_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n393_), .A2(new_n394_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n397_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(new_n207_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  OR3_X1    g206(.A1(new_n399_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n399_), .B2(new_n403_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n394_), .A2(KEYINPUT29), .ZN(new_n411_));
  XOR2_X1   g210(.A(G211gat), .B(G218gat), .Z(new_n412_));
  INV_X1    g211(.A(G204gat), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n413_), .A2(G197gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(G197gat), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n417_));
  AOI21_X1  g216(.A(new_n412_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT90), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n414_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n415_), .A2(new_n419_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT21), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT21), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n416_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n412_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G233gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n411_), .A2(new_n428_), .A3(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n435_), .B(KEYINPUT92), .Z(new_n436_));
  XOR2_X1   g235(.A(G78gat), .B(G106gat), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n428_), .A2(KEYINPUT93), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n418_), .A2(new_n423_), .B1(new_n426_), .B2(new_n412_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT93), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n411_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n433_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n436_), .A2(new_n438_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n394_), .A2(KEYINPUT29), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT28), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G22gat), .B(G50gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n438_), .B1(new_n436_), .B2(new_n445_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n447_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n454_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n456_), .B2(new_n446_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n410_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G183gat), .A2(G190gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT23), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(G183gat), .B2(G190gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT22), .B(G169gat), .ZN(new_n462_));
  INV_X1    g261(.A(G176gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G169gat), .A2(G176gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n465_), .B(KEYINPUT95), .Z(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT96), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n461_), .A2(KEYINPUT96), .A3(new_n464_), .A4(new_n466_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(G169gat), .A2(G176gat), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n472_), .A2(KEYINPUT24), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n460_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT25), .B(G183gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT26), .B(G190gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(KEYINPUT24), .A3(new_n465_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n480_), .A2(KEYINPUT94), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(KEYINPUT94), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n475_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n428_), .B1(new_n471_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT22), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(G169gat), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n463_), .B(new_n488_), .C1(new_n462_), .C2(new_n486_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n461_), .A2(new_n465_), .A3(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n478_), .A2(new_n460_), .A3(new_n473_), .A4(new_n479_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n485_), .B1(new_n493_), .B2(new_n440_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n484_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G226gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT19), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n471_), .A2(new_n483_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n440_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n497_), .ZN(new_n501_));
  OAI211_X1 g300(.A(KEYINPUT20), .B(new_n501_), .C1(new_n493_), .C2(new_n440_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G8gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT18), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G64gat), .B(G92gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n498_), .A2(new_n504_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n502_), .B1(new_n440_), .B2(new_n499_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n501_), .B1(new_n484_), .B2(new_n494_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n508_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n513_), .A3(KEYINPUT97), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT97), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n515_), .B(new_n508_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT27), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n514_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n495_), .A2(new_n497_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n483_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n520_), .A2(new_n467_), .A3(new_n439_), .A4(new_n442_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n428_), .B2(new_n492_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n501_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n508_), .B1(new_n519_), .B2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(KEYINPUT27), .A3(new_n510_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n518_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n458_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n514_), .A2(new_n516_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT33), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT98), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n409_), .B(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n407_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT99), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n400_), .A2(new_n397_), .A3(new_n402_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n529_), .A2(new_n532_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT100), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT100), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n529_), .A2(new_n532_), .A3(new_n539_), .A4(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n509_), .A2(KEYINPUT32), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n511_), .A2(new_n512_), .A3(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n410_), .A2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n519_), .B2(new_n524_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT102), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n538_), .A2(new_n540_), .A3(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n455_), .A2(new_n457_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n528_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n492_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(G99gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n492_), .B(KEYINPUT30), .ZN(new_n554_));
  INV_X1    g353(.A(G99gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT85), .B(G43gat), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G227gat), .A2(G233gat), .ZN(new_n561_));
  INV_X1    g360(.A(G15gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(G71gat), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n553_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n560_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n566_), .A2(KEYINPUT87), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n564_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n565_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n558_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n567_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n566_), .A3(KEYINPUT87), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n568_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n393_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(new_n576_), .A3(new_n393_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT103), .B1(new_n550_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n579_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(new_n577_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT103), .ZN(new_n584_));
  INV_X1    g383(.A(new_n549_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n537_), .A2(KEYINPUT100), .B1(new_n544_), .B2(new_n546_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n586_), .B2(new_n540_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n583_), .B(new_n584_), .C1(new_n587_), .C2(new_n528_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n581_), .A2(new_n588_), .ZN(new_n589_));
  AOI211_X1 g388(.A(new_n527_), .B(new_n585_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n410_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n296_), .A2(new_n297_), .A3(new_n250_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n250_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n297_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n294_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n249_), .B(new_n246_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n255_), .A2(new_n297_), .A3(new_n296_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n593_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G169gat), .B(G197gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n604_), .B(new_n605_), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(KEYINPUT82), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT82), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n597_), .A2(new_n602_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT83), .Z(new_n612_));
  NAND3_X1  g411(.A1(new_n592_), .A2(KEYINPUT104), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT104), .B1(new_n592_), .B2(new_n612_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n322_), .B(new_n370_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n616_), .A2(G1gat), .A3(new_n410_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n581_), .A2(new_n588_), .B1(new_n590_), .B2(new_n410_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n284_), .A2(new_n271_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n611_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n369_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT105), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n321_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n623_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n410_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n619_), .A2(new_n620_), .A3(new_n629_), .ZN(G1324gat));
  NAND3_X1  g429(.A1(new_n623_), .A2(new_n527_), .A3(new_n627_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n631_), .A2(new_n632_), .A3(G8gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n631_), .B2(G8gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n527_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n635_), .A2(new_n289_), .ZN(new_n636_));
  OAI22_X1  g435(.A1(new_n633_), .A2(new_n634_), .B1(new_n616_), .B2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1325gat));
  OAI21_X1  g438(.A(G15gat), .B1(new_n628_), .B2(new_n583_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT41), .Z(new_n641_));
  NAND2_X1  g440(.A1(new_n580_), .A2(new_n562_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n616_), .B2(new_n642_), .ZN(G1326gat));
  OAI21_X1  g442(.A(G22gat), .B1(new_n628_), .B2(new_n549_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT42), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n549_), .A2(G22gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n616_), .B2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(new_n321_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n622_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n370_), .B(new_n650_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n651_), .A2(G29gat), .A3(new_n410_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT108), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n589_), .A2(new_n653_), .A3(new_n591_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n653_), .A2(KEYINPUT43), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n654_), .B(new_n287_), .C1(new_n621_), .C2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT107), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT43), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(KEYINPUT43), .ZN(new_n659_));
  INV_X1    g458(.A(new_n287_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n621_), .B2(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n656_), .A2(new_n658_), .A3(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n626_), .A2(new_n648_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(KEYINPUT44), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n410_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n656_), .A2(new_n658_), .A3(new_n661_), .A4(new_n663_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n665_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n652_), .B1(new_n669_), .B2(G29gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT109), .ZN(G1328gat));
  INV_X1    g470(.A(new_n651_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT110), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n635_), .A2(G36gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n674_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT110), .B1(new_n651_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n664_), .A2(new_n668_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G36gat), .B1(new_n681_), .B2(new_n635_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n675_), .A2(new_n677_), .A3(KEYINPUT45), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n680_), .A2(new_n682_), .A3(KEYINPUT46), .A4(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1329gat));
  INV_X1    g487(.A(G43gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n651_), .B2(new_n583_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n664_), .A2(G43gat), .A3(new_n580_), .A4(new_n668_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT47), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n692_), .A2(new_n696_), .A3(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1330gat));
  INV_X1    g497(.A(G50gat), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n681_), .A2(new_n699_), .A3(new_n549_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G50gat), .B1(new_n672_), .B2(new_n585_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1331gat));
  NAND2_X1  g501(.A1(new_n369_), .A2(new_n624_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n621_), .A2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(new_n322_), .ZN(new_n705_));
  INV_X1    g504(.A(G57gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n665_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n321_), .A2(new_n612_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n623_), .A2(new_n369_), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n410_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1332gat));
  OAI21_X1  g510(.A(G64gat), .B1(new_n709_), .B2(new_n635_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT48), .ZN(new_n713_));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n705_), .A2(new_n714_), .A3(new_n527_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT112), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n709_), .B2(new_n583_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n705_), .A2(new_n721_), .A3(new_n580_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1334gat));
  OAI21_X1  g522(.A(G78gat), .B1(new_n709_), .B2(new_n549_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n549_), .A2(G78gat), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT114), .Z(new_n727_));
  NAND2_X1  g526(.A1(new_n705_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n648_), .A2(new_n703_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT115), .Z(new_n731_));
  NAND4_X1  g530(.A1(new_n656_), .A2(new_n731_), .A3(new_n658_), .A4(new_n661_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT116), .ZN(new_n733_));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n410_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n704_), .A2(new_n650_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n207_), .A3(new_n665_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(G1336gat));
  OAI21_X1  g537(.A(G92gat), .B1(new_n733_), .B2(new_n635_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n208_), .A3(new_n527_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1337gat));
  NOR2_X1   g540(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n662_), .A2(new_n580_), .A3(new_n731_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G99gat), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n736_), .A2(new_n203_), .A3(new_n205_), .A4(new_n580_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n742_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n746_), .B(new_n747_), .Z(G1338gat));
  NAND3_X1  g547(.A1(new_n736_), .A2(new_n204_), .A3(new_n585_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n732_), .A2(new_n549_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n204_), .B1(new_n751_), .B2(KEYINPUT118), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT118), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n732_), .B2(new_n549_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n750_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n662_), .A2(KEYINPUT118), .A3(new_n585_), .A4(new_n731_), .ZN(new_n756_));
  AND4_X1   g555(.A1(new_n750_), .A2(new_n756_), .A3(G106gat), .A4(new_n754_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n749_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n749_), .C1(new_n755_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n590_), .A2(new_n665_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n595_), .A2(new_n596_), .A3(new_n594_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n593_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n606_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n607_), .B1(new_n597_), .B2(new_n602_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT120), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n603_), .A2(new_n606_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT120), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n765_), .A2(new_n606_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n769_), .B(new_n770_), .C1(new_n771_), .C2(new_n764_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n364_), .A2(new_n768_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n345_), .A2(new_n774_), .A3(new_n348_), .ZN(new_n775_));
  AND4_X1   g574(.A1(new_n333_), .A2(new_n337_), .A3(new_n338_), .A4(new_n342_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n333_), .A2(new_n337_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(KEYINPUT55), .B1(new_n777_), .B2(new_n349_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n360_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n360_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(KEYINPUT119), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT119), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n779_), .A2(new_n785_), .A3(KEYINPUT56), .A4(new_n360_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n611_), .A2(new_n363_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n773_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT121), .B1(new_n789_), .B2(new_n622_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n786_), .A2(new_n787_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n360_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n781_), .B(new_n359_), .C1(new_n775_), .C2(new_n778_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n792_), .B1(new_n795_), .B2(KEYINPUT119), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n791_), .B(new_n649_), .C1(new_n796_), .C2(new_n773_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n790_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT122), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n790_), .A2(new_n797_), .A3(KEYINPUT122), .A4(new_n798_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n789_), .A2(new_n798_), .A3(new_n622_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n772_), .A2(new_n768_), .A3(new_n363_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n794_), .B2(new_n793_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n804_), .B(KEYINPUT58), .C1(new_n794_), .C2(new_n793_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n287_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n803_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n801_), .A2(new_n802_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n321_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n708_), .A2(new_n660_), .A3(new_n370_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n813_), .A2(KEYINPUT54), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(KEYINPUT54), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n763_), .B1(new_n812_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(G113gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n611_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n814_), .A2(new_n815_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n321_), .B2(new_n811_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n821_), .B2(new_n763_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n763_), .A2(KEYINPUT59), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n648_), .B1(new_n810_), .B2(new_n799_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n826_), .A2(new_n612_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n819_), .B1(new_n827_), .B2(new_n818_), .ZN(G1340gat));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n369_), .B(new_n825_), .C1(new_n817_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT60), .B1(new_n369_), .B2(new_n833_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n821_), .A2(new_n763_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n822_), .A2(KEYINPUT123), .A3(new_n369_), .A4(new_n825_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n832_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G120gat), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT124), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n836_), .A2(KEYINPUT60), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n835_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n833_), .B1(new_n844_), .B2(new_n837_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT124), .B1(new_n845_), .B2(new_n841_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(G1341gat));
  INV_X1    g646(.A(G127gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n817_), .A2(new_n848_), .A3(new_n648_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n826_), .A2(new_n648_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n848_), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n817_), .A2(new_n852_), .A3(new_n622_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n826_), .A2(new_n287_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n852_), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n812_), .A2(new_n816_), .ZN(new_n856_));
  NOR4_X1   g655(.A1(new_n580_), .A2(new_n527_), .A3(new_n410_), .A4(new_n549_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n624_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(new_n375_), .ZN(G1344gat));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n370_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n376_), .ZN(G1345gat));
  NOR2_X1   g661(.A1(new_n858_), .A2(new_n321_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT61), .B(G155gat), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  OAI21_X1  g664(.A(G162gat), .B1(new_n858_), .B2(new_n660_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n649_), .A2(G162gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n858_), .B2(new_n867_), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n820_), .A2(new_n824_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n585_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n583_), .A2(new_n635_), .A3(new_n665_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G169gat), .B1(new_n872_), .B2(new_n624_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n874_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n870_), .A2(new_n462_), .A3(new_n611_), .A4(new_n871_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(G1348gat));
  OAI21_X1  g677(.A(new_n463_), .B1(new_n872_), .B2(new_n370_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n821_), .A2(new_n585_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n880_), .A2(G176gat), .A3(new_n369_), .A4(new_n871_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1349gat));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n648_), .A3(new_n871_), .ZN(new_n883_));
  INV_X1    g682(.A(G183gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n871_), .A2(new_n648_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n476_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n883_), .A2(new_n884_), .B1(new_n870_), .B2(new_n886_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n872_), .B2(new_n660_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n622_), .A2(new_n477_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n872_), .B2(new_n889_), .ZN(G1351gat));
  NOR3_X1   g689(.A1(new_n580_), .A2(new_n665_), .A3(new_n549_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT126), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n635_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n856_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n611_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g696(.A1(new_n894_), .A2(new_n370_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n413_), .ZN(G1353gat));
  XNOR2_X1  g698(.A(KEYINPUT63), .B(G211gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n895_), .A2(new_n648_), .A3(new_n900_), .ZN(new_n901_));
  OAI22_X1  g700(.A1(new_n894_), .A2(new_n321_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT127), .Z(G1354gat));
  OAI21_X1  g703(.A(G218gat), .B1(new_n894_), .B2(new_n660_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n649_), .A2(G218gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n894_), .B2(new_n906_), .ZN(G1355gat));
endmodule


