//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n208_), .B(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G229gat), .A2(G233gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n213_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n208_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n213_), .B2(new_n208_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n216_), .B1(new_n220_), .B2(new_n215_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G113gat), .B(G141gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G169gat), .B(G197gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n221_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT96), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT85), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G141gat), .A2(G148gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT87), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT1), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n234_), .B(new_n235_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n233_), .B(KEYINPUT3), .Z(new_n242_));
  XOR2_X1   g041(.A(new_n235_), .B(KEYINPUT2), .Z(new_n243_));
  OAI211_X1 g042(.A(new_n237_), .B(new_n239_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n232_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n241_), .A2(new_n230_), .A3(new_n244_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n250_), .B2(new_n247_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT91), .Z(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n252_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G1gat), .B(G29gat), .ZN(new_n257_));
  INV_X1    g056(.A(G85gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G57gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n254_), .A2(new_n255_), .A3(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(G197gat), .B(G204gat), .Z(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(KEYINPUT21), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(KEYINPUT21), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n245_), .B2(KEYINPUT29), .ZN(new_n271_));
  AND2_X1   g070(.A1(G228gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G78gat), .B(G106gat), .Z(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n273_), .A2(new_n274_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n276_), .B2(KEYINPUT88), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT89), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n245_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT28), .B(G22gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(G50gat), .B1(new_n245_), .B2(KEYINPUT29), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n280_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n273_), .A2(new_n274_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT88), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n277_), .A2(new_n278_), .A3(new_n284_), .A4(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n273_), .A2(new_n274_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n273_), .A2(KEYINPUT88), .A3(new_n274_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n287_), .A2(new_n289_), .A3(new_n284_), .A4(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT89), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  OAI22_X1  g092(.A1(new_n276_), .A2(new_n275_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n265_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT20), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT23), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(G183gat), .A3(G190gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n300_), .A2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT90), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT24), .ZN(new_n309_));
  OR3_X1    g108(.A1(new_n305_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n307_), .B(KEYINPUT81), .Z(new_n311_));
  INV_X1    g110(.A(KEYINPUT24), .ZN(new_n312_));
  AND2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT25), .B(G183gat), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n306_), .B1(new_n305_), .B2(new_n309_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n310_), .A2(new_n314_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT22), .B(G169gat), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n313_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(new_n301_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n270_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n296_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G226gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT19), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT26), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n315_), .A2(KEYINPUT79), .B1(KEYINPUT80), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G183gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(KEYINPUT25), .ZN(new_n336_));
  OAI221_X1 g135(.A(new_n334_), .B1(KEYINPUT79), .B2(new_n336_), .C1(KEYINPUT80), .C2(new_n317_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n301_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n311_), .A2(new_n312_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n314_), .A4(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n323_), .B1(new_n305_), .B2(new_n324_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n270_), .A3(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n328_), .A2(new_n331_), .A3(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n320_), .A2(new_n270_), .A3(new_n325_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT20), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT93), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n341_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n327_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT93), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n349_), .A3(KEYINPUT20), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n343_), .B1(new_n351_), .B2(new_n330_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G92gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT18), .B(G64gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  OR2_X1    g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n344_), .A2(new_n348_), .A3(KEYINPUT20), .A4(new_n331_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n328_), .A2(new_n342_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n358_), .B(new_n356_), .C1(new_n359_), .C2(new_n331_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(KEYINPUT27), .A3(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT94), .B(KEYINPUT27), .ZN(new_n362_));
  INV_X1    g161(.A(new_n356_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n331_), .B1(new_n328_), .B2(new_n342_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n358_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n360_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT95), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n368_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n295_), .B(new_n361_), .C1(new_n369_), .C2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n356_), .A2(KEYINPUT32), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n358_), .B(new_n373_), .C1(new_n359_), .C2(new_n331_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n265_), .B(new_n374_), .C1(new_n352_), .C2(new_n373_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n261_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT92), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n251_), .A2(new_n252_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT33), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n378_), .A2(new_n379_), .B1(new_n264_), .B2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n264_), .A2(new_n380_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n375_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n293_), .A2(new_n294_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n372_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n347_), .B(KEYINPUT30), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT84), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT31), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT83), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G15gat), .B(G43gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n394_), .B(new_n395_), .Z(new_n396_));
  NAND3_X1  g195(.A1(new_n389_), .A2(new_n390_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n390_), .B1(new_n389_), .B2(new_n396_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT86), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n397_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n388_), .A2(KEYINPUT84), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(new_n232_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n400_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n227_), .B1(new_n387_), .B2(new_n409_), .ZN(new_n410_));
  AOI211_X1 g209(.A(KEYINPUT96), .B(new_n408_), .C1(new_n372_), .C2(new_n386_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n409_), .A2(new_n265_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n361_), .B1(new_n371_), .B2(new_n369_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n385_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n226_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT37), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G190gat), .B(G218gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G134gat), .B(G162gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n422_), .A2(KEYINPUT36), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G232gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT34), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT67), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT66), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G99gat), .A2(G106gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT66), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n431_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT7), .ZN(new_n440_));
  INV_X1    g239(.A(G99gat), .ZN(new_n441_));
  INV_X1    g240(.A(G106gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT67), .A3(new_n427_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n430_), .A2(new_n434_), .A3(new_n439_), .A4(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G85gat), .B(G92gat), .Z(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT68), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(new_n449_), .A3(new_n446_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(KEYINPUT8), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT69), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n432_), .A2(new_n433_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n443_), .A3(new_n427_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT8), .B1(new_n455_), .B2(KEYINPUT65), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n456_), .B(new_n446_), .C1(KEYINPUT65), .C2(new_n455_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n448_), .A2(KEYINPUT69), .A3(KEYINPUT8), .A4(new_n450_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n213_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT10), .B(G99gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT64), .B(G106gat), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n446_), .A2(KEYINPUT9), .ZN(new_n465_));
  INV_X1    g264(.A(G92gat), .ZN(new_n466_));
  OR3_X1    g265(.A1(new_n258_), .A2(new_n466_), .A3(KEYINPUT9), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .A4(new_n454_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n459_), .A2(new_n460_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n218_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(new_n459_), .B2(new_n468_), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT35), .B(new_n425_), .C1(new_n470_), .C2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n472_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n425_), .A2(KEYINPUT35), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n425_), .A2(KEYINPUT35), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .A4(new_n469_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n423_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT72), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n422_), .A2(KEYINPUT36), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n477_), .A3(new_n423_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT73), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n418_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n478_), .A2(new_n480_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n479_), .B1(new_n484_), .B2(new_n418_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n482_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n459_), .A2(new_n468_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G57gat), .B(G64gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT70), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT11), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G71gat), .B(G78gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT11), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n492_), .A2(new_n497_), .A3(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n490_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n459_), .A2(new_n468_), .A3(new_n499_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G230gat), .A2(G233gat), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n490_), .A2(KEYINPUT12), .A3(new_n500_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n503_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n504_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n505_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G120gat), .B(G148gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G204gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT5), .B(G176gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n516_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n508_), .A2(new_n511_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT13), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(KEYINPUT13), .A3(new_n519_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n489_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G231gat), .A2(G233gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT74), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n208_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n499_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G183gat), .B(G211gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G127gat), .B(G155gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n529_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n534_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(KEYINPUT17), .B2(new_n538_), .ZN(new_n539_));
  AND4_X1   g338(.A1(KEYINPUT76), .A2(new_n529_), .A3(KEYINPUT17), .A4(new_n538_), .ZN(new_n540_));
  AOI21_X1  g339(.A(KEYINPUT76), .B1(new_n529_), .B2(new_n536_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT77), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n525_), .A2(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT78), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT78), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n417_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(new_n203_), .A3(new_n265_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT38), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT97), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n387_), .A2(new_n409_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT96), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n387_), .A2(new_n409_), .A3(new_n227_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n416_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n524_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n225_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n479_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT98), .B1(new_n483_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT98), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n542_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n555_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n203_), .B1(new_n566_), .B2(new_n265_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n548_), .B1(new_n549_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n551_), .A2(new_n568_), .ZN(G1324gat));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n547_), .A2(new_n570_), .A3(new_n204_), .A4(new_n414_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n417_), .A2(new_n204_), .A3(new_n546_), .A4(new_n545_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT99), .B1(new_n572_), .B2(new_n415_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT40), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n555_), .A2(new_n564_), .A3(new_n414_), .A4(new_n565_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(G8gat), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n576_), .B2(G8gat), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n574_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n575_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n582_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n574_), .A2(new_n580_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT40), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n584_), .B1(new_n588_), .B2(new_n581_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n586_), .A2(new_n589_), .ZN(G1325gat));
  INV_X1    g389(.A(G15gat), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n566_), .B2(new_n408_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT41), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n547_), .A2(new_n591_), .A3(new_n408_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(G1326gat));
  INV_X1    g394(.A(G22gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n385_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n566_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT103), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT42), .Z(new_n600_));
  NAND3_X1  g399(.A1(new_n547_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1327gat));
  INV_X1    g401(.A(new_n563_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n557_), .A2(new_n543_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(G29gat), .B1(new_n606_), .B2(new_n265_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n265_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n555_), .A2(new_n489_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT43), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT43), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n555_), .A2(new_n611_), .A3(new_n489_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n605_), .B(KEYINPUT104), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT44), .ZN(new_n617_));
  INV_X1    g416(.A(new_n614_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT105), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n617_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n608_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n607_), .B1(new_n622_), .B2(G29gat), .ZN(G1328gat));
  XNOR2_X1  g422(.A(new_n414_), .B(KEYINPUT106), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n555_), .A2(new_n563_), .A3(new_n605_), .A4(new_n624_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n625_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT107), .B1(new_n625_), .B2(G36gat), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n626_), .A2(KEYINPUT45), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT45), .B1(new_n626_), .B2(new_n627_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n415_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n631_));
  INV_X1    g430(.A(G36gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT46), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n630_), .B(KEYINPUT46), .C1(new_n631_), .C2(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1329gat));
  INV_X1    g436(.A(KEYINPUT47), .ZN(new_n638_));
  INV_X1    g437(.A(G43gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n616_), .A2(new_n621_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(new_n408_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n606_), .A2(new_n639_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n409_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n638_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n409_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n645_));
  OAI221_X1 g444(.A(KEYINPUT47), .B1(new_n409_), .B2(new_n642_), .C1(new_n645_), .C2(new_n639_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1330gat));
  AOI21_X1  g446(.A(KEYINPUT44), .B1(new_n615_), .B2(KEYINPUT105), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n619_), .A2(new_n620_), .A3(new_n617_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n597_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n640_), .A2(KEYINPUT108), .A3(new_n597_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(G50gat), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(G50gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n606_), .A2(new_n655_), .A3(new_n597_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1331gat));
  AOI21_X1  g456(.A(new_n556_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n489_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n543_), .A2(new_n226_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n658_), .A2(new_n659_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G57gat), .B1(new_n662_), .B2(new_n265_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(new_n603_), .A3(new_n661_), .ZN(new_n664_));
  INV_X1    g463(.A(G57gat), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(new_n608_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n663_), .A2(new_n666_), .ZN(G1332gat));
  INV_X1    g466(.A(new_n624_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G64gat), .B1(new_n664_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT48), .ZN(new_n670_));
  INV_X1    g469(.A(G64gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n662_), .A2(new_n671_), .A3(new_n624_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1333gat));
  OAI21_X1  g472(.A(G71gat), .B1(new_n664_), .B2(new_n409_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT49), .ZN(new_n675_));
  INV_X1    g474(.A(new_n662_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n409_), .A2(G71gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT109), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n676_), .B2(new_n678_), .ZN(G1334gat));
  OAI21_X1  g478(.A(G78gat), .B1(new_n664_), .B2(new_n385_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n385_), .A2(G78gat), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT111), .Z(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n676_), .B2(new_n684_), .ZN(G1335gat));
  NOR3_X1   g484(.A1(new_n556_), .A2(new_n225_), .A3(new_n543_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n604_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G85gat), .B1(new_n688_), .B2(new_n265_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n613_), .A2(new_n686_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT112), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n613_), .A2(KEYINPUT112), .A3(new_n686_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n608_), .A2(new_n258_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n689_), .B1(new_n694_), .B2(new_n695_), .ZN(G1336gat));
  AOI21_X1  g495(.A(G92gat), .B1(new_n688_), .B2(new_n414_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n668_), .A2(new_n466_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n694_), .B2(new_n698_), .ZN(G1337gat));
  NAND3_X1  g498(.A1(new_n692_), .A2(new_n408_), .A3(new_n693_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G99gat), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n687_), .A2(new_n461_), .A3(new_n409_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT113), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT51), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(new_n703_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1338gat));
  NAND3_X1  g507(.A1(new_n688_), .A2(new_n463_), .A3(new_n597_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n613_), .A2(new_n597_), .A3(new_n686_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT52), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(G106gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G106gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g514(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n659_), .A2(new_n556_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT77), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n542_), .B(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(KEYINPUT114), .A3(new_n225_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT114), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n543_), .B2(new_n226_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n717_), .B1(new_n718_), .B2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n525_), .B(new_n716_), .C1(new_n723_), .C2(new_n721_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT118), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n519_), .A2(KEYINPUT116), .A3(new_n225_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT116), .B1(new_n519_), .B2(new_n225_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n503_), .A2(new_n504_), .A3(new_n507_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n510_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n508_), .A2(new_n734_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n503_), .A2(new_n506_), .A3(KEYINPUT55), .A4(new_n507_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n733_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n516_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT56), .B1(new_n737_), .B2(new_n516_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n731_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n221_), .A2(new_n224_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n214_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(new_n215_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n220_), .B(KEYINPUT117), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n215_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n741_), .B1(new_n745_), .B2(new_n224_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n520_), .A2(new_n746_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n740_), .A2(new_n747_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n728_), .B1(new_n748_), .B2(KEYINPUT57), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT57), .ZN(new_n750_));
  INV_X1    g549(.A(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n737_), .A2(new_n516_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n516_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n751_), .B1(new_n756_), .B2(new_n731_), .ZN(new_n757_));
  OAI211_X1 g556(.A(KEYINPUT118), .B(new_n750_), .C1(new_n757_), .C2(new_n563_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n748_), .A2(KEYINPUT57), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n519_), .B(new_n746_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n756_), .A2(KEYINPUT58), .A3(new_n519_), .A4(new_n746_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n489_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n749_), .A2(new_n758_), .A3(new_n759_), .A4(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n727_), .B1(new_n765_), .B2(new_n542_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n608_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n409_), .A2(new_n597_), .A3(new_n414_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G113gat), .B1(new_n770_), .B2(new_n225_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n759_), .A2(new_n764_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n748_), .A2(KEYINPUT57), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n720_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n727_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n768_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n776_), .A2(KEYINPUT59), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n265_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n769_), .A2(KEYINPUT59), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n225_), .A2(G113gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n771_), .B1(new_n781_), .B2(new_n782_), .ZN(G1340gat));
  NAND3_X1  g582(.A1(new_n779_), .A2(new_n780_), .A3(new_n524_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT60), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n556_), .A2(G120gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n769_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G120gat), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1341gat));
  AOI21_X1  g589(.A(G127gat), .B1(new_n770_), .B2(new_n543_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n565_), .A2(G127gat), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n791_), .B1(new_n781_), .B2(new_n793_), .ZN(G1342gat));
  AOI21_X1  g593(.A(G134gat), .B1(new_n770_), .B2(new_n563_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n489_), .A2(G134gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n781_), .B2(new_n796_), .ZN(G1343gat));
  NOR3_X1   g596(.A1(new_n624_), .A2(new_n385_), .A3(new_n408_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n767_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n225_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g601(.A1(new_n799_), .A2(new_n556_), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT119), .B(G148gat), .Z(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(G1345gat));
  OR3_X1    g604(.A1(new_n799_), .A2(G155gat), .A3(new_n720_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n807_));
  OAI21_X1  g606(.A(G155gat), .B1(new_n799_), .B2(new_n720_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1346gat));
  AND3_X1   g610(.A1(new_n800_), .A2(G162gat), .A3(new_n489_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G162gat), .B1(new_n800_), .B2(new_n563_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1347gat));
  NAND2_X1  g613(.A1(new_n624_), .A2(new_n413_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT121), .ZN(new_n816_));
  OR3_X1    g615(.A1(new_n776_), .A2(new_n597_), .A3(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(G169gat), .B1(new_n817_), .B2(new_n226_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n776_), .A2(new_n597_), .A3(new_n816_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(new_n225_), .A3(new_n321_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  MUX2_X1   g620(.A(new_n818_), .B(new_n821_), .S(KEYINPUT62), .Z(G1348gat));
  NOR2_X1   g621(.A1(new_n766_), .A2(new_n597_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n816_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(G176gat), .A3(new_n524_), .A4(new_n824_), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(KEYINPUT122), .Z(new_n826_));
  AOI21_X1  g625(.A(G176gat), .B1(new_n819_), .B2(new_n524_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(G1349gat));
  NAND3_X1  g627(.A1(new_n823_), .A2(new_n543_), .A3(new_n824_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n565_), .A2(new_n315_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n829_), .A2(new_n335_), .B1(new_n819_), .B2(new_n831_), .ZN(G1350gat));
  OAI21_X1  g631(.A(G190gat), .B1(new_n817_), .B2(new_n659_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n819_), .A2(new_n563_), .A3(new_n317_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(G1351gat));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n765_), .A2(new_n542_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n775_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n624_), .A2(new_n409_), .A3(new_n295_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n836_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n766_), .A2(KEYINPUT123), .A3(new_n839_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n225_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT125), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n838_), .A2(new_n836_), .A3(new_n840_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT123), .B1(new_n766_), .B2(new_n839_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n226_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT125), .B1(new_n849_), .B2(KEYINPUT124), .ZN(new_n850_));
  AOI21_X1  g649(.A(G197gat), .B1(new_n849_), .B2(KEYINPUT124), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n846_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n846_), .B2(new_n850_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1352gat));
  NOR2_X1   g653(.A1(new_n841_), .A2(new_n842_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n556_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n857_));
  AND2_X1   g656(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n856_), .B2(new_n857_), .ZN(G1353gat));
  INV_X1    g659(.A(new_n855_), .ZN(new_n861_));
  AOI211_X1 g660(.A(KEYINPUT63), .B(G211gat), .C1(new_n861_), .C2(new_n565_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT63), .B(G211gat), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n855_), .A2(new_n542_), .A3(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1354gat));
  AOI21_X1  g664(.A(G218gat), .B1(new_n861_), .B2(new_n563_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n855_), .A2(new_n659_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(G218gat), .ZN(G1355gat));
endmodule


