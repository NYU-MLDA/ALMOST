//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT71), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(KEYINPUT71), .A2(G183gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT75), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n218_), .A2(KEYINPUT75), .A3(G183gat), .A4(G190gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT74), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n217_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G169gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n213_), .A2(KEYINPUT25), .A3(new_n214_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT72), .A3(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n237_), .A2(G183gat), .B1(new_n216_), .B2(KEYINPUT26), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT72), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(new_n216_), .B2(KEYINPUT26), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n234_), .A2(new_n236_), .A3(new_n238_), .A4(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT73), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n225_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n224_), .A2(KEYINPUT73), .A3(KEYINPUT23), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n219_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT24), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(G169gat), .B2(G176gat), .ZN(new_n248_));
  INV_X1    g047(.A(G169gat), .ZN(new_n249_));
  INV_X1    g048(.A(G176gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n246_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n241_), .A2(new_n245_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n233_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT88), .ZN(new_n256_));
  XOR2_X1   g055(.A(G211gat), .B(G218gat), .Z(new_n257_));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT87), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n262_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n264_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n263_), .A2(KEYINPUT87), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n261_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT86), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(KEYINPUT86), .A3(new_n261_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n256_), .B(new_n265_), .C1(new_n269_), .C2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n262_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n256_), .B1(new_n278_), .B2(new_n265_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n255_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT20), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n245_), .B1(G183gat), .B2(G190gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT96), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n232_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n224_), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT74), .B1(new_n224_), .B2(KEYINPUT23), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n221_), .A2(new_n222_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n246_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT94), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT25), .B(G183gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n251_), .B1(new_n248_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT24), .B1(new_n249_), .B2(new_n250_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT93), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n295_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n292_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n246_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(KEYINPUT94), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n302_), .A2(KEYINPUT95), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT95), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n300_), .B1(new_n303_), .B2(KEYINPUT94), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n290_), .A2(new_n291_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT94), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n306_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n285_), .B1(new_n305_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n265_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n281_), .B1(new_n314_), .B2(KEYINPUT97), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT97), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n316_), .A3(new_n313_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n210_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(KEYINPUT88), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(new_n275_), .A3(new_n254_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(KEYINPUT20), .A3(new_n210_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n265_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n274_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n323_), .B2(new_n277_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT95), .B1(new_n302_), .B2(new_n304_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n307_), .A2(new_n310_), .A3(new_n306_), .ZN(new_n326_));
  AOI22_X1  g125(.A1(new_n325_), .A2(new_n326_), .B1(new_n232_), .B2(new_n284_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n321_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n206_), .B1(new_n318_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n330_), .A2(KEYINPUT78), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(KEYINPUT78), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G113gat), .B(G120gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n331_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n339_));
  INV_X1    g138(.A(G141gat), .ZN(new_n340_));
  INV_X1    g139(.A(G148gat), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .A4(KEYINPUT82), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT82), .ZN(new_n343_));
  OAI22_X1  g142(.A1(new_n343_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n342_), .A2(new_n344_), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G155gat), .ZN(new_n350_));
  INV_X1    g149(.A(G162gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(KEYINPUT81), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(G155gat), .B2(G162gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n349_), .A2(new_n352_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(KEYINPUT1), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(G155gat), .A3(G162gat), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n357_), .A2(new_n352_), .A3(new_n354_), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n340_), .A2(new_n341_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n345_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n338_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n336_), .A2(new_n337_), .A3(new_n362_), .A4(new_n356_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n338_), .A2(new_n367_), .A3(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n364_), .A2(new_n371_), .A3(new_n365_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n372_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n377_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n370_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n371_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT33), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(KEYINPUT33), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n379_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT97), .B1(new_n327_), .B2(new_n324_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n280_), .A2(KEYINPUT20), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n317_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n328_), .B1(new_n389_), .B2(new_n209_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n205_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n329_), .A2(new_n386_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT98), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n369_), .A2(new_n371_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n382_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n377_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(KEYINPUT99), .A3(new_n383_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT99), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(new_n380_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n285_), .B(new_n324_), .C1(new_n304_), .C2(new_n302_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(KEYINPUT20), .A3(new_n320_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n209_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n389_), .B2(new_n209_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n401_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n390_), .A2(new_n406_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n329_), .A2(new_n386_), .A3(new_n391_), .A4(KEYINPUT98), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n394_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415_));
  INV_X1    g214(.A(new_n232_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n290_), .B2(new_n217_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n241_), .A2(new_n245_), .A3(new_n252_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n415_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT76), .B(G43gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT77), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n288_), .A2(new_n289_), .B1(new_n216_), .B2(new_n215_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n253_), .B(KEYINPUT30), .C1(new_n423_), .C2(new_n416_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n419_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427_));
  INV_X1    g226(.A(G15gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G71gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G99gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n425_), .A2(new_n426_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT30), .B1(new_n233_), .B2(new_n253_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n424_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n421_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n419_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n431_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n414_), .B1(new_n433_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n432_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n431_), .A3(new_n437_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT79), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n338_), .B(KEYINPUT31), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT79), .A4(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n413_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(KEYINPUT80), .A3(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT29), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n356_), .A2(new_n362_), .A3(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G22gat), .B(G50gat), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT83), .B(KEYINPUT28), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n453_), .A2(new_n454_), .ZN(new_n459_));
  OR3_X1    g258(.A1(new_n456_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n452_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT84), .B(G228gat), .ZN(new_n464_));
  INV_X1    g263(.A(G233gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT85), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n319_), .A2(new_n468_), .A3(new_n275_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n324_), .B2(new_n463_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G78gat), .B(G106gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n471_), .B(KEYINPUT89), .Z(new_n472_));
  AND3_X1   g271(.A1(new_n469_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n462_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT90), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n462_), .B(KEYINPUT90), .C1(new_n473_), .C2(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n469_), .A2(new_n470_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n462_), .B1(new_n480_), .B2(new_n471_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n473_), .A2(KEYINPUT91), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n473_), .A2(KEYINPUT91), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n451_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n401_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n449_), .A2(KEYINPUT80), .A3(new_n446_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT80), .B1(new_n449_), .B2(new_n446_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n485_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n444_), .A2(new_n447_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(new_n484_), .A3(new_n479_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n489_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT27), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n390_), .A2(new_n205_), .ZN(new_n497_));
  AOI211_X1 g296(.A(new_n206_), .B(new_n328_), .C1(new_n389_), .C2(new_n209_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n405_), .A2(new_n206_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n391_), .A3(KEYINPUT27), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n412_), .A2(new_n488_), .B1(new_n495_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G29gat), .B(G36gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n505_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT15), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  INV_X1    g309(.A(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G8gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n508_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(new_n516_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n518_), .B(new_n516_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT70), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n529_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n521_), .A2(new_n524_), .A3(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n503_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G230gat), .A2(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G85gat), .B(G92gat), .Z(new_n537_));
  NAND2_X1  g336(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT7), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n539_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT65), .B(G92gat), .Z(new_n548_));
  INV_X1    g347(.A(G85gat), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(KEYINPUT9), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n544_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n537_), .A2(KEYINPUT9), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT64), .ZN(new_n553_));
  XOR2_X1   g352(.A(KEYINPUT10), .B(G99gat), .Z(new_n554_));
  INV_X1    g353(.A(G106gat), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n554_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n551_), .B(new_n552_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n558_));
  OAI221_X1 g357(.A(new_n539_), .B1(KEYINPUT66), .B2(KEYINPUT8), .C1(new_n544_), .C2(new_n541_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n547_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n563_));
  XOR2_X1   g362(.A(G71gat), .B(G78gat), .Z(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n560_), .A2(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n547_), .A2(new_n558_), .A3(new_n559_), .A4(new_n567_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(KEYINPUT12), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT12), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n560_), .A2(new_n572_), .A3(new_n568_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n536_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n535_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G120gat), .B(G148gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n581_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n583_), .B(new_n584_), .C1(KEYINPUT68), .C2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n567_), .B(new_n516_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595_));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT16), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  OR3_X1    g398(.A1(new_n594_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(KEYINPUT17), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n594_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n560_), .A2(new_n518_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT69), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT34), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT35), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n604_), .A2(new_n605_), .A3(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n608_), .A2(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n604_), .A2(new_n610_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n560_), .A2(new_n509_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(KEYINPUT36), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n611_), .B(new_n612_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n620_), .B(KEYINPUT36), .Z(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n617_), .B2(new_n622_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT37), .B1(new_n624_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n617_), .A2(new_n622_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n629_), .B(new_n623_), .C1(new_n630_), .C2(new_n626_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n534_), .A2(new_n590_), .A3(new_n603_), .A4(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT101), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n633_), .B(KEYINPUT100), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n636_), .A2(new_n639_), .A3(new_n511_), .A4(new_n489_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n624_), .A2(new_n627_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n503_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n590_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n603_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n533_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n401_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n640_), .A2(new_n641_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n642_), .A2(new_n649_), .A3(new_n650_), .ZN(G1324gat));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n652_));
  INV_X1    g451(.A(new_n648_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n499_), .A2(new_n501_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(KEYINPUT102), .A3(G8gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n512_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(KEYINPUT102), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT103), .B(new_n652_), .C1(new_n657_), .C2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n502_), .A2(G8gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n636_), .A2(new_n639_), .A3(new_n661_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n658_), .A2(KEYINPUT102), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n656_), .A3(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n662_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n660_), .A2(new_n662_), .A3(KEYINPUT40), .A4(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n648_), .B2(new_n451_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT41), .Z(new_n672_));
  INV_X1    g471(.A(new_n451_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n635_), .A2(new_n428_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1326gat));
  OAI21_X1  g474(.A(G22gat), .B1(new_n648_), .B2(new_n486_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT42), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n486_), .A2(G22gat), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT104), .Z(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n637_), .B2(new_n679_), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n646_), .A2(new_n643_), .ZN(new_n681_));
  NOR4_X1   g480(.A1(new_n503_), .A2(new_n533_), .A3(new_n645_), .A4(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n489_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n503_), .B2(new_n632_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(new_n632_), .ZN(new_n686_));
  AND4_X1   g485(.A1(new_n484_), .A2(new_n479_), .A3(new_n446_), .A4(new_n449_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n451_), .B2(new_n485_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n688_), .A2(new_n654_), .A3(new_n489_), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n392_), .A2(new_n393_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n487_), .B1(new_n690_), .B2(new_n411_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n685_), .B(new_n686_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n684_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n533_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n646_), .A2(new_n694_), .A3(new_n590_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT44), .B1(new_n693_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  AOI211_X1 g497(.A(new_n698_), .B(new_n695_), .C1(new_n684_), .C2(new_n692_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n489_), .A2(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n683_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT46), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n697_), .A2(new_n699_), .A3(new_n502_), .ZN(new_n706_));
  INV_X1    g505(.A(G36gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n693_), .A2(new_n696_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n698_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n696_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n654_), .A3(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n708_), .A2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n502_), .A2(G36gat), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n682_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n682_), .B2(new_n716_), .ZN(new_n718_));
  OAI22_X1  g517(.A1(new_n717_), .A2(new_n718_), .B1(new_n703_), .B2(KEYINPUT46), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n704_), .B1(new_n714_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n704_), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n722_), .B(new_n719_), .C1(new_n708_), .C2(new_n713_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1329gat));
  AOI21_X1  g523(.A(G43gat), .B1(new_n682_), .B2(new_n673_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n493_), .A2(G43gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n700_), .B2(new_n726_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n682_), .B2(new_n485_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n485_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n700_), .B2(new_n730_), .ZN(G1331gat));
  NOR2_X1   g530(.A1(new_n503_), .A2(new_n694_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n686_), .A2(new_n590_), .A3(new_n646_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n401_), .B1(new_n734_), .B2(KEYINPUT108), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(KEYINPUT108), .B2(new_n734_), .ZN(new_n736_));
  INV_X1    g535(.A(G57gat), .ZN(new_n737_));
  AND4_X1   g536(.A1(new_n533_), .A2(new_n644_), .A3(new_n645_), .A4(new_n603_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n489_), .B2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n739_), .B2(new_n737_), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n736_), .A2(new_n737_), .B1(new_n738_), .B2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n738_), .B2(new_n654_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n734_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n743_), .A3(new_n654_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n738_), .B2(new_n673_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT49), .Z(new_n752_));
  NAND3_X1  g551(.A1(new_n747_), .A2(new_n750_), .A3(new_n673_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1334gat));
  INV_X1    g553(.A(G78gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n738_), .B2(new_n485_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT50), .Z(new_n757_));
  NAND2_X1  g556(.A1(new_n485_), .A2(new_n755_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT111), .Z(new_n759_));
  OAI21_X1  g558(.A(new_n757_), .B1(new_n734_), .B2(new_n759_), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n603_), .A2(new_n694_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n693_), .A2(new_n645_), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n401_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n681_), .A2(new_n590_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n732_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n549_), .A3(new_n489_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n763_), .A2(new_n767_), .ZN(G1336gat));
  AOI21_X1  g567(.A(G92gat), .B1(new_n766_), .B2(new_n654_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n762_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n654_), .A2(new_n548_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n770_), .B2(new_n771_), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n762_), .B2(new_n451_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n493_), .A2(new_n554_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n765_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g575(.A1(new_n693_), .A2(new_n485_), .A3(new_n645_), .A4(new_n761_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n777_), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT113), .B1(new_n777_), .B2(G106gat), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n780_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n765_), .A2(G106gat), .A3(new_n486_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  OR3_X1    g586(.A1(new_n781_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n781_), .B2(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1339gat));
  INV_X1    g589(.A(G113gat), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n694_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n792_), .B2(new_n791_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n654_), .A2(new_n401_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n574_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n571_), .A2(new_n536_), .A3(new_n573_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n582_), .B1(new_n574_), .B2(new_n799_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n517_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n522_), .A2(new_n520_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .A4(new_n529_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n532_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n529_), .A3(new_n809_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(KEYINPUT117), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n583_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n803_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT118), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n806_), .B(new_n815_), .C1(new_n817_), .C2(new_n804_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n814_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(KEYINPUT58), .C1(new_n804_), .C2(new_n817_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n686_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n801_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n824_), .A2(new_n574_), .A3(new_n799_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n574_), .A2(new_n799_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n581_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n825_), .A2(new_n827_), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n828_));
  NOR2_X1   g627(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n802_), .A2(new_n803_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n533_), .B1(new_n576_), .B2(new_n582_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n828_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n832_), .A2(new_n833_), .B1(new_n585_), .B2(new_n813_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n828_), .A2(new_n831_), .A3(new_n830_), .A4(KEYINPUT116), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n643_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n823_), .B1(new_n836_), .B2(KEYINPUT57), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n832_), .A2(new_n833_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n585_), .A2(new_n813_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n835_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n643_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n646_), .B1(new_n837_), .B2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n632_), .A2(new_n533_), .A3(new_n590_), .A4(new_n603_), .ZN(new_n846_));
  XOR2_X1   g645(.A(new_n846_), .B(KEYINPUT54), .Z(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n798_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT59), .B1(new_n849_), .B2(new_n687_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n632_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n842_), .A2(new_n843_), .B1(new_n851_), .B2(new_n822_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n836_), .A2(KEYINPUT57), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n603_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n687_), .B(new_n797_), .C1(new_n854_), .C2(new_n847_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n796_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n849_), .A2(KEYINPUT59), .A3(new_n687_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n856_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(KEYINPUT119), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n795_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n855_), .ZN(new_n863_));
  AOI21_X1  g662(.A(G113gat), .B1(new_n863_), .B2(new_n694_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT121), .B1(new_n862_), .B2(new_n864_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n859_), .A2(new_n860_), .A3(KEYINPUT119), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT119), .B1(new_n859_), .B2(new_n860_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n794_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  INV_X1    g668(.A(new_n864_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n865_), .A2(new_n871_), .ZN(G1340gat));
  AOI21_X1  g671(.A(new_n590_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(KEYINPUT122), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n590_), .A2(G120gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n863_), .B1(KEYINPUT60), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n873_), .B2(KEYINPUT122), .ZN(new_n877_));
  OAI21_X1  g676(.A(G120gat), .B1(new_n874_), .B2(new_n877_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n876_), .A2(KEYINPUT60), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1341gat));
  INV_X1    g679(.A(G127gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n863_), .A2(new_n881_), .A3(new_n603_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n646_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1342gat));
  INV_X1    g683(.A(G134gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n863_), .A2(new_n885_), .A3(new_n643_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n632_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1343gat));
  NAND3_X1  g687(.A1(new_n849_), .A2(new_n485_), .A3(new_n451_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n533_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT123), .B(G141gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n590_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n341_), .ZN(G1345gat));
  NOR2_X1   g693(.A1(new_n889_), .A2(new_n646_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT61), .B(G155gat), .Z(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n889_), .B2(new_n632_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n643_), .A2(new_n351_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n889_), .B2(new_n899_), .ZN(G1347gat));
  NAND2_X1  g699(.A1(new_n845_), .A2(new_n848_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n502_), .A2(new_n489_), .A3(new_n485_), .A4(new_n451_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n249_), .B1(new_n903_), .B2(new_n694_), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT62), .Z(new_n905_));
  INV_X1    g704(.A(new_n903_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT22), .B(G169gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n694_), .A2(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT124), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n905_), .B1(new_n906_), .B2(new_n909_), .ZN(G1348gat));
  NAND2_X1  g709(.A1(new_n903_), .A2(new_n645_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g711(.A1(new_n903_), .A2(new_n603_), .ZN(new_n913_));
  OR3_X1    g712(.A1(new_n913_), .A2(KEYINPUT125), .A3(new_n293_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT125), .B1(new_n913_), .B2(new_n293_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n215_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n906_), .B2(new_n632_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n903_), .A2(new_n294_), .A3(new_n643_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1351gat));
  NOR3_X1   g719(.A1(new_n502_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n901_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n533_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT126), .B(G197gat), .Z(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1352gat));
  INV_X1    g724(.A(new_n922_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n645_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g727(.A1(new_n922_), .A2(new_n646_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  AND2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n932_), .B1(new_n929_), .B2(new_n930_), .ZN(G1354gat));
  AND3_X1   g732(.A1(new_n926_), .A2(G218gat), .A3(new_n686_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n922_), .A2(new_n841_), .ZN(new_n935_));
  OR2_X1    g734(.A1(new_n935_), .A2(KEYINPUT127), .ZN(new_n936_));
  AOI21_X1  g735(.A(G218gat), .B1(new_n935_), .B2(KEYINPUT127), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n934_), .B1(new_n936_), .B2(new_n937_), .ZN(G1355gat));
endmodule


