//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_;
  INV_X1    g000(.A(G197gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT89), .B1(new_n202_), .B2(G204gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT89), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(G197gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n202_), .A2(G204gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n209_));
  OR2_X1    g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n205_), .A2(G197gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(new_n207_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n211_), .B1(KEYINPUT21), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n210_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT91), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n210_), .A2(KEYINPUT91), .A3(new_n214_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n211_), .A2(KEYINPUT21), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n208_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT86), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  INV_X1    g030(.A(G141gat), .ZN(new_n232_));
  INV_X1    g031(.A(G148gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(new_n231_), .A3(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(KEYINPUT2), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n237_));
  OR4_X1    g036(.A1(new_n237_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n237_), .B2(KEYINPUT3), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n222_), .B1(new_n223_), .B2(new_n242_), .ZN(new_n243_));
  AND3_X1   g042(.A1(KEYINPUT92), .A2(G228gat), .A3(G233gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT92), .B1(G228gat), .B2(G233gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n245_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G22gat), .B(G50gat), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n235_), .A2(new_n241_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT28), .B1(new_n251_), .B2(KEYINPUT29), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n251_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n253_), .A2(KEYINPUT88), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT88), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n257_), .B2(new_n252_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n250_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT88), .B1(new_n253_), .B2(new_n254_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n257_), .A2(new_n256_), .A3(new_n252_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n250_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n264_), .A2(KEYINPUT93), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n259_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n249_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G15gat), .B(G43gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT31), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G227gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(KEYINPUT83), .B(KEYINPUT23), .Z(new_n275_));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(KEYINPUT23), .B2(new_n276_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT81), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT84), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT84), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n278_), .A2(new_n285_), .A3(new_n282_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n279_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT24), .A3(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(KEYINPUT82), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT25), .B(G183gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G190gat), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n290_), .A2(KEYINPUT82), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n284_), .A2(new_n286_), .A3(new_n291_), .A4(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n276_), .A2(KEYINPUT23), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G176gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT22), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT85), .B1(new_n302_), .B2(G169gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT22), .B(G169gat), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n301_), .B(new_n303_), .C1(new_n304_), .C2(KEYINPUT85), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(new_n289_), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n295_), .A2(KEYINPUT30), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT30), .B1(new_n295_), .B2(new_n306_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n274_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G127gat), .B(G134gat), .Z(new_n311_));
  XOR2_X1   g110(.A(G113gat), .B(G120gat), .Z(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n295_), .A2(new_n306_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT30), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n274_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n307_), .A3(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n310_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n314_), .B1(new_n310_), .B2(new_n319_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n271_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n308_), .A2(new_n309_), .A3(new_n274_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n318_), .B1(new_n317_), .B2(new_n307_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n313_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n270_), .A3(new_n320_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n264_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n262_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n249_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n259_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n268_), .A2(new_n323_), .A3(new_n327_), .A4(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G8gat), .B(G36gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT18), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G64gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G92gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n340_), .A2(KEYINPUT32), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT97), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n292_), .B(KEYINPUT94), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n293_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n290_), .A2(new_n297_), .A3(new_n282_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n304_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n289_), .B1(new_n349_), .B2(G176gat), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(new_n278_), .B2(new_n299_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n343_), .B1(new_n222_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n315_), .B2(new_n222_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT19), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n315_), .A2(new_n222_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n217_), .A2(new_n218_), .B1(new_n208_), .B2(new_n220_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n351_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n343_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n357_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n342_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n242_), .A2(new_n314_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n251_), .A2(new_n313_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(KEYINPUT4), .A3(new_n369_), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n242_), .A2(KEYINPUT4), .A3(new_n314_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT95), .Z(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G1gat), .B(G29gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT0), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G57gat), .ZN(new_n379_));
  INV_X1    g178(.A(G85gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n376_), .A2(KEYINPUT98), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n376_), .A2(new_n382_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n374_), .A2(new_n375_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT98), .B1(new_n385_), .B2(new_n381_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n359_), .A2(new_n362_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n357_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n357_), .B2(new_n355_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n341_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n367_), .A2(new_n383_), .A3(new_n387_), .A4(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT96), .Z(new_n394_));
  NAND2_X1  g193(.A1(new_n368_), .A2(new_n369_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n382_), .B1(new_n396_), .B2(new_n373_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n394_), .A2(new_n397_), .B1(new_n398_), .B2(new_n384_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n358_), .A2(new_n340_), .A3(new_n364_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n365_), .A2(new_n339_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n376_), .A2(KEYINPUT33), .A3(new_n382_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n335_), .B1(new_n392_), .B2(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n387_), .A2(KEYINPUT99), .A3(new_n383_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT99), .B1(new_n387_), .B2(new_n383_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n332_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n327_), .B(new_n323_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n327_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n270_), .B1(new_n326_), .B2(new_n320_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n268_), .B(new_n334_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n407_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n401_), .A2(new_n400_), .ZN(new_n415_));
  XOR2_X1   g214(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n400_), .A2(KEYINPUT100), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n390_), .A2(new_n339_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT100), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n358_), .A2(new_n420_), .A3(new_n340_), .A4(new_n364_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT27), .A4(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n404_), .B1(new_n414_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G230gat), .ZN(new_n425_));
  INV_X1    g224(.A(G233gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT11), .ZN(new_n428_));
  INV_X1    g227(.A(G64gat), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n429_), .A2(G57gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(G57gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G57gat), .B(G64gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT11), .ZN(new_n434_));
  INV_X1    g233(.A(G71gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT68), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT68), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G71gat), .ZN(new_n438_));
  INV_X1    g237(.A(G78gat), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n432_), .B(new_n434_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n440_), .A2(new_n441_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n443_), .B2(new_n434_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT7), .ZN(new_n446_));
  INV_X1    g245(.A(G99gat), .ZN(new_n447_));
  INV_X1    g246(.A(G106gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT8), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n455_));
  NAND2_X1  g254(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n455_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n448_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(G85gat), .B2(G92gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G92gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n380_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n463_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n462_), .B1(new_n467_), .B2(KEYINPUT9), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n453_), .B1(new_n459_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT66), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n380_), .A2(new_n463_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n449_), .A2(KEYINPUT8), .A3(new_n451_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(new_n474_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n450_), .A2(KEYINPUT67), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  OAI221_X1 g282(.A(new_n479_), .B1(KEYINPUT67), .B2(new_n450_), .C1(new_n480_), .C2(new_n474_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n445_), .B1(new_n476_), .B2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n485_), .B(new_n444_), .C1(new_n469_), .C2(new_n475_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT12), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n454_), .A2(new_n456_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT64), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n492_));
  AOI21_X1  g291(.A(G106gat), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n466_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(G92gat), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT9), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n461_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n452_), .B1(new_n493_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n475_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n485_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT12), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n445_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n427_), .B1(new_n489_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n427_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G120gat), .B(G148gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(new_n205_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT5), .B(G176gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  OR3_X1    g313(.A1(new_n505_), .A2(new_n507_), .A3(new_n513_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT13), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(KEYINPUT13), .A3(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G169gat), .B(G197gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G141gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT80), .B(G113gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  XNOR2_X1  g323(.A(G29gat), .B(G36gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G43gat), .B(G50gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(G8gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT74), .B(G22gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G15gat), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT75), .B(G1gat), .Z(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n533_), .B2(G8gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(G1gat), .B1(new_n531_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n531_), .A2(G1gat), .A3(new_n534_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n529_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(G8gat), .A3(new_n535_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n528_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT15), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n527_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n538_), .A2(new_n540_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT79), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n538_), .A2(new_n540_), .A3(new_n528_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n547_), .B1(new_n542_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n524_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n524_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n542_), .A2(new_n552_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n550_), .B(new_n555_), .C1(new_n556_), .C2(new_n547_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n520_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n424_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT69), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT34), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n499_), .A2(new_n500_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n527_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n544_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT35), .B(new_n565_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n545_), .A2(new_n502_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .A4(new_n567_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT70), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G190gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(G218gat), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n578_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT36), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n575_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(KEYINPUT36), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n570_), .A2(new_n587_), .A3(new_n574_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT71), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n570_), .A2(new_n587_), .A3(KEYINPUT71), .A4(new_n574_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n586_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT37), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT72), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n590_), .A2(KEYINPUT72), .A3(new_n591_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT73), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n585_), .B(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n596_), .B(new_n597_), .C1(new_n575_), .C2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n594_), .B1(new_n600_), .B2(KEYINPUT37), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT78), .ZN(new_n603_));
  XOR2_X1   g402(.A(G183gat), .B(G211gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT17), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n607_), .A2(KEYINPUT17), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n538_), .A2(new_n540_), .A3(new_n444_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT76), .Z(new_n614_));
  AOI21_X1  g413(.A(new_n444_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n612_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n614_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n615_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n618_), .B2(new_n611_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n609_), .B(new_n610_), .C1(new_n616_), .C2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n616_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(new_n608_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n601_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n562_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n407_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n533_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n629_), .A2(KEYINPUT38), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(KEYINPUT38), .ZN(new_n631_));
  INV_X1    g430(.A(new_n593_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n424_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n561_), .A2(new_n624_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n627_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n630_), .A2(new_n631_), .A3(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  OAI21_X1  g437(.A(G8gat), .B1(new_n635_), .B2(new_n423_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n423_), .A2(G8gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n562_), .A2(new_n625_), .A3(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT102), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n646_));
  AND2_X1   g445(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n647_));
  OR3_X1    g446(.A1(new_n639_), .A2(new_n640_), .A3(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n645_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n646_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n638_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n645_), .A2(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT104), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n645_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(KEYINPUT40), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n655_), .ZN(G1325gat));
  NOR2_X1   g455(.A1(new_n411_), .A2(new_n412_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G15gat), .B1(new_n635_), .B2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT41), .Z(new_n659_));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n657_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n626_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n662_), .ZN(G1326gat));
  NOR2_X1   g462(.A1(new_n408_), .A2(new_n409_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G22gat), .B1(new_n635_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  INV_X1    g465(.A(G22gat), .ZN(new_n667_));
  INV_X1    g466(.A(new_n664_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n626_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(G1327gat));
  NAND2_X1  g469(.A1(new_n410_), .A2(new_n413_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n627_), .A3(new_n423_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n404_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n624_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n561_), .A2(new_n675_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n674_), .A2(new_n632_), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n407_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n601_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n424_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n674_), .A2(new_n681_), .A3(new_n601_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n676_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n683_), .A2(KEYINPUT44), .A3(new_n676_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n407_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n678_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  INV_X1    g489(.A(new_n423_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n686_), .A2(new_n691_), .A3(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT105), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n686_), .A2(new_n694_), .A3(new_n691_), .A4(new_n687_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n693_), .A2(G36gat), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n677_), .A2(new_n697_), .A3(new_n691_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT45), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n696_), .A2(KEYINPUT46), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  NOR2_X1   g503(.A1(new_n657_), .A2(G43gat), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n677_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n688_), .A2(new_n661_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G43gat), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT47), .B(new_n706_), .C1(new_n707_), .C2(G43gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n677_), .B2(new_n668_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n668_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n688_), .B2(new_n714_), .ZN(G1331gat));
  AND4_X1   g514(.A1(new_n623_), .A2(new_n620_), .A3(new_n554_), .A4(new_n557_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n520_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n633_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n627_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n520_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(new_n558_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n674_), .A2(new_n625_), .A3(new_n721_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n627_), .A2(G57gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(new_n722_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n429_), .A3(new_n691_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G64gat), .B1(new_n718_), .B2(new_n423_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(KEYINPUT48), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(KEYINPUT48), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT106), .Z(G1333gat));
  OAI21_X1  g530(.A(G71gat), .B1(new_n718_), .B2(new_n657_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT49), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n657_), .A2(G71gat), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT107), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n722_), .B2(new_n735_), .ZN(G1334gat));
  OAI21_X1  g535(.A(G78gat), .B1(new_n718_), .B2(new_n664_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT50), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n725_), .A2(new_n439_), .A3(new_n668_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT108), .ZN(G1335gat));
  NAND2_X1  g540(.A1(new_n721_), .A2(new_n624_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n683_), .A2(new_n743_), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n627_), .B(new_n744_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n424_), .A2(new_n742_), .A3(new_n593_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n407_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT109), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1336gat));
  OAI21_X1  g548(.A(G92gat), .B1(new_n744_), .B2(new_n423_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(new_n463_), .A3(new_n691_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1337gat));
  OAI21_X1  g551(.A(G99gat), .B1(new_n744_), .B2(new_n657_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n746_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n661_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n746_), .A2(new_n448_), .A3(new_n668_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n424_), .A2(KEYINPUT43), .A3(new_n679_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n681_), .B1(new_n674_), .B2(new_n601_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n668_), .B(new_n743_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(G106gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G106gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n758_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT110), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n758_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n766_), .A2(KEYINPUT53), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT53), .B1(new_n766_), .B2(new_n768_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1339gat));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT114), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n558_), .A2(new_n515_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n427_), .A2(KEYINPUT112), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n488_), .A2(KEYINPUT12), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n444_), .B1(new_n501_), .B2(new_n485_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n566_), .A2(KEYINPUT12), .A3(new_n444_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT55), .B(new_n776_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(KEYINPUT55), .B2(new_n505_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n489_), .A2(new_n504_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n776_), .B1(new_n783_), .B2(KEYINPUT55), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n775_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT55), .B1(new_n779_), .B2(new_n780_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(KEYINPUT112), .A3(new_n427_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n506_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n787_), .A2(new_n790_), .A3(KEYINPUT113), .A4(new_n781_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n513_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n791_), .A4(new_n513_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n774_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n542_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n524_), .B(new_n797_), .C1(new_n556_), .C2(new_n548_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n516_), .A2(new_n557_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n593_), .B(new_n773_), .C1(new_n796_), .C2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n557_), .A2(new_n798_), .A3(new_n515_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n601_), .B1(new_n803_), .B2(KEYINPUT58), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n805_), .B(new_n802_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n801_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n774_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n787_), .A2(new_n781_), .A3(new_n790_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n512_), .B1(new_n809_), .B2(new_n775_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n791_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n795_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n799_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n773_), .B1(new_n814_), .B2(new_n593_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n624_), .B1(new_n807_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n716_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n716_), .A2(KEYINPUT111), .A3(new_n518_), .A4(new_n519_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n679_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT54), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n679_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n816_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n691_), .A2(new_n627_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n413_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT115), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT116), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n827_), .A2(new_n834_), .A3(new_n831_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n558_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n832_), .A2(KEYINPUT59), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n827_), .A2(new_n840_), .A3(new_n831_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(new_n558_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n843_), .B2(new_n837_), .ZN(G1340gat));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n520_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n720_), .B2(G120gat), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n833_), .A2(new_n835_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G120gat), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1341gat));
  AOI21_X1  g650(.A(G127gat), .B1(new_n836_), .B2(new_n675_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n675_), .A2(G127gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT117), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n842_), .B2(new_n854_), .ZN(G1342gat));
  NAND3_X1  g654(.A1(new_n833_), .A2(new_n632_), .A3(new_n835_), .ZN(new_n856_));
  INV_X1    g655(.A(G134gat), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT118), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n856_), .A2(new_n860_), .A3(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n601_), .A2(G134gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT119), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n859_), .A2(new_n861_), .B1(new_n842_), .B2(new_n863_), .ZN(G1343gat));
  AOI21_X1  g663(.A(new_n410_), .B1(new_n816_), .B2(new_n826_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n828_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n559_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n232_), .ZN(G1344gat));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n720_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n233_), .ZN(G1345gat));
  NOR2_X1   g669(.A1(new_n866_), .A2(new_n624_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT61), .B(G155gat), .Z(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  OAI21_X1  g672(.A(G162gat), .B1(new_n866_), .B2(new_n679_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n593_), .A2(G162gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n866_), .B2(new_n875_), .ZN(G1347gat));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n423_), .A2(new_n407_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n829_), .ZN(new_n879_));
  AOI211_X1 g678(.A(new_n559_), .B(new_n879_), .C1(new_n816_), .C2(new_n826_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G169gat), .B1(new_n880_), .B2(KEYINPUT120), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n816_), .B2(new_n826_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n882_), .A2(KEYINPUT120), .A3(new_n558_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n877_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885_));
  INV_X1    g684(.A(new_n879_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n827_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n887_), .B2(new_n559_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n880_), .A2(KEYINPUT120), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n880_), .A2(new_n304_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n884_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n884_), .A2(KEYINPUT121), .A3(new_n890_), .A4(new_n891_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1348gat));
  NAND2_X1  g695(.A1(new_n882_), .A2(new_n520_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g697(.A1(new_n882_), .A2(new_n675_), .A3(new_n344_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n900_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G183gat), .B1(new_n882_), .B2(new_n675_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n887_), .B2(new_n679_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT123), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n882_), .A2(new_n632_), .A3(new_n293_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1351gat));
  NAND2_X1  g707(.A1(new_n865_), .A2(new_n878_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n558_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n911_), .A2(KEYINPUT124), .A3(new_n202_), .ZN(new_n912_));
  AOI21_X1  g711(.A(KEYINPUT124), .B1(new_n911_), .B2(new_n202_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n911_), .A2(new_n202_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n910_), .A2(new_n520_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n205_), .A2(KEYINPUT125), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1353gat));
  NOR2_X1   g717(.A1(new_n909_), .A2(new_n624_), .ZN(new_n919_));
  OR2_X1    g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT127), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  OR3_X1    g720(.A1(new_n919_), .A2(KEYINPUT127), .A3(new_n920_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT63), .B(G211gat), .Z(new_n923_));
  NAND2_X1  g722(.A1(new_n919_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n919_), .A2(KEYINPUT126), .A3(new_n923_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n921_), .A2(new_n922_), .B1(new_n926_), .B2(new_n927_), .ZN(G1354gat));
  OAI21_X1  g727(.A(G218gat), .B1(new_n909_), .B2(new_n679_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n632_), .A2(new_n582_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n909_), .B2(new_n930_), .ZN(G1355gat));
endmodule


