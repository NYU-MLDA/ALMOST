//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n969_, new_n970_, new_n971_, new_n972_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G43gat), .B(G50gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n210_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n206_), .A2(new_n207_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n209_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n216_), .B(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n217_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(new_n208_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n218_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n215_), .B(new_n213_), .C1(new_n221_), .C2(new_n208_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n218_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(KEYINPUT77), .A3(new_n218_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n226_), .B1(new_n225_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G113gat), .B(G141gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT78), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G169gat), .B(G197gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n233_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT100), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT83), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n247_), .A3(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(KEYINPUT23), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT81), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(KEYINPUT24), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n254_), .B1(G169gat), .B2(G176gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT26), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G190gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT79), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT25), .B(G183gat), .ZN(new_n260_));
  INV_X1    g059(.A(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT26), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT80), .B1(new_n259_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n258_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n262_), .A4(new_n260_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n250_), .A2(new_n256_), .A3(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n244_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT84), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(new_n241_), .B2(KEYINPUT23), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n271_), .B(new_n273_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n274_));
  INV_X1    g073(.A(G183gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n261_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n278_));
  INV_X1    g077(.A(G169gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n270_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n284_), .A2(new_n288_), .A3(new_n285_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n240_), .B1(new_n283_), .B2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n293_));
  NAND2_X1  g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n280_), .B1(new_n250_), .B2(new_n276_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n255_), .A2(KEYINPUT98), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n255_), .A2(KEYINPUT98), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n252_), .A3(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n262_), .A2(new_n258_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n300_), .A2(new_n260_), .B1(new_n254_), .B2(new_n251_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n274_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n296_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n295_), .B1(new_n304_), .B2(new_n291_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n270_), .A2(new_n282_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n289_), .A2(new_n290_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(KEYINPUT100), .A3(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n292_), .A2(new_n305_), .A3(KEYINPUT20), .A4(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n307_), .B1(new_n296_), .B2(new_n303_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n270_), .A2(new_n282_), .A3(new_n291_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(KEYINPUT20), .A3(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n312_), .A2(KEYINPUT99), .A3(new_n295_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT99), .B1(new_n312_), .B2(new_n295_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G8gat), .B(G36gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT18), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n319_), .B(new_n309_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT27), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n312_), .A2(new_n295_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT104), .B1(new_n296_), .B2(new_n303_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT104), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n245_), .A2(KEYINPUT83), .B1(KEYINPUT23), .B2(new_n241_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n329_), .A2(new_n248_), .B1(new_n275_), .B2(new_n261_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n328_), .B(new_n302_), .C1(new_n330_), .C2(new_n280_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n291_), .A3(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n292_), .A2(new_n332_), .A3(KEYINPUT20), .A4(new_n308_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n326_), .B1(new_n333_), .B2(new_n295_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n322_), .B(KEYINPUT27), .C1(new_n319_), .C2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT92), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT91), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT91), .B1(new_n343_), .B2(KEYINPUT92), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n342_), .A2(new_n343_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT2), .Z(new_n347_));
  OAI211_X1 g146(.A(new_n337_), .B(new_n338_), .C1(new_n345_), .C2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n336_), .B1(KEYINPUT1), .B2(new_n338_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(KEYINPUT1), .B2(new_n338_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n340_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n346_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n348_), .A2(new_n352_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT28), .B1(new_n357_), .B2(KEYINPUT29), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G22gat), .B(G50gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n356_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(KEYINPUT96), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT96), .ZN(new_n365_));
  INV_X1    g164(.A(new_n363_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n360_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n307_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n369_));
  INV_X1    g168(.A(G233gat), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n370_), .A2(KEYINPUT93), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(KEYINPUT93), .ZN(new_n372_));
  OAI21_X1  g171(.A(G228gat), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT94), .B1(new_n369_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n291_), .B1(new_n357_), .B2(KEYINPUT29), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT94), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n373_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT95), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n369_), .A2(new_n380_), .A3(new_n374_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT95), .B1(new_n376_), .B2(new_n373_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G78gat), .B(G106gat), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n379_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n364_), .B(new_n368_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n379_), .A2(new_n383_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n384_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n364_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n386_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n325_), .A2(new_n335_), .A3(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n306_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT87), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT86), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G15gat), .B(G43gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n283_), .A2(new_n396_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n270_), .A2(new_n282_), .A3(new_n396_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n398_), .A2(new_n405_), .A3(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n397_), .A2(KEYINPUT87), .A3(new_n404_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT90), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G127gat), .B(G134gat), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n414_), .A2(KEYINPUT88), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(KEYINPUT88), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G113gat), .B(G120gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n415_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT90), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n410_), .A2(new_n426_), .A3(new_n411_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n413_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  AOI211_X1 g227(.A(new_n426_), .B(new_n425_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n353_), .A2(new_n422_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n357_), .A2(new_n421_), .A3(new_n420_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(KEYINPUT4), .A3(new_n432_), .ZN(new_n433_));
  OR3_X1    g232(.A1(new_n353_), .A2(new_n422_), .A3(KEYINPUT4), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT101), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n431_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G85gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n444_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n437_), .A2(new_n438_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n428_), .A2(new_n430_), .A3(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n395_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n424_), .B1(new_n412_), .B2(KEYINPUT90), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n429_), .B1(new_n452_), .B2(new_n427_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(KEYINPUT33), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n437_), .A2(new_n455_), .A3(new_n438_), .A4(new_n446_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n431_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n444_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT103), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT103), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n457_), .A2(new_n461_), .A3(new_n444_), .A4(new_n458_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n454_), .A2(new_n456_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n319_), .A2(KEYINPUT32), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n309_), .B(new_n465_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n466_), .B(new_n448_), .C1(new_n334_), .C2(new_n465_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n394_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n387_), .A2(new_n364_), .A3(new_n388_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n368_), .A2(new_n364_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(new_n391_), .B2(new_n386_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n470_), .A2(new_n472_), .A3(new_n448_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n325_), .A2(new_n473_), .A3(new_n335_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n453_), .B1(new_n469_), .B2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n451_), .B1(new_n475_), .B2(KEYINPUT105), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT105), .ZN(new_n477_));
  INV_X1    g276(.A(new_n335_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT27), .B1(new_n321_), .B2(new_n322_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n389_), .A2(new_n449_), .A3(new_n393_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n470_), .A2(new_n472_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n482_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n477_), .B1(new_n484_), .B2(new_n453_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n239_), .B1(new_n476_), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G190gat), .B(G218gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT75), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G134gat), .B(G162gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n490_), .A2(new_n491_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G232gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT35), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT73), .Z(new_n498_));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT10), .B(G99gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n503_), .B1(new_n504_), .B2(G106gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT64), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT9), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT9), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT64), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(KEYINPUT9), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n507_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  AOI211_X1 g319(.A(KEYINPUT65), .B(new_n518_), .C1(new_n512_), .C2(new_n515_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n506_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n500_), .A2(new_n502_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n526_));
  INV_X1    g325(.A(G99gat), .ZN(new_n527_));
  INV_X1    g326(.A(G106gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(KEYINPUT66), .B(new_n515_), .C1(new_n525_), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT67), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n534_), .B(new_n515_), .C1(new_n525_), .C2(new_n531_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(KEYINPUT8), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n532_), .A2(KEYINPUT67), .A3(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT68), .B(new_n506_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n524_), .A2(new_n536_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n216_), .B(KEYINPUT15), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n498_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n496_), .A2(KEYINPUT35), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G85gat), .B(G92gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n530_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n547_), .B2(new_n503_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n534_), .B1(new_n548_), .B2(KEYINPUT66), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n535_), .A2(KEYINPUT8), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n538_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n519_), .B1(new_n544_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT65), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n516_), .A2(new_n507_), .A3(new_n519_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n505_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n543_), .B1(new_n557_), .B2(new_n216_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n542_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT76), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT76), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n542_), .A2(new_n561_), .A3(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n498_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n536_), .A2(new_n216_), .A3(new_n538_), .A4(new_n522_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n565_), .B1(KEYINPUT35), .B2(new_n496_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n540_), .A2(new_n541_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(KEYINPUT74), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n556_), .B(new_n523_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n551_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n220_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT74), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n564_), .B1(new_n568_), .B2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n492_), .B(new_n493_), .C1(new_n563_), .C2(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n542_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n561_), .B1(new_n542_), .B2(new_n558_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n558_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n567_), .A2(KEYINPUT74), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n498_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n578_), .A2(new_n581_), .A3(new_n491_), .A4(new_n490_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n575_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n575_), .A2(new_n582_), .A3(KEYINPUT37), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G57gat), .B(G64gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT11), .ZN(new_n590_));
  XOR2_X1   g389(.A(G71gat), .B(G78gat), .Z(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n589_), .A2(KEYINPUT11), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n590_), .A2(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n222_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601_));
  XOR2_X1   g400(.A(G127gat), .B(G155gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n600_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(KEYINPUT17), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n600_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n588_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n594_), .A2(KEYINPUT12), .A3(new_n595_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n540_), .A2(new_n613_), .B1(new_n557_), .B2(new_n596_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n596_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n551_), .B2(new_n556_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(new_n615_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n557_), .A2(new_n596_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n617_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n615_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT5), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n626_), .B(new_n627_), .Z(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n620_), .A2(new_n624_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT70), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n629_), .B1(new_n620_), .B2(new_n624_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n620_), .A2(new_n624_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n628_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT70), .B1(new_n636_), .B2(new_n630_), .ZN(new_n637_));
  OAI22_X1  g436(.A1(new_n634_), .A2(new_n637_), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n632_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n636_), .A2(KEYINPUT70), .A3(new_n630_), .ZN(new_n640_));
  XOR2_X1   g439(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n611_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n486_), .A2(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(G1gat), .A3(new_n449_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n645_), .A2(new_n609_), .A3(new_n239_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n453_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT105), .B(new_n652_), .C1(new_n481_), .C2(new_n483_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n395_), .A2(new_n450_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n469_), .A2(new_n474_), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT105), .B1(new_n656_), .B2(new_n652_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n583_), .B(new_n651_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n476_), .A2(new_n485_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n661_), .A2(KEYINPUT107), .A3(new_n583_), .A4(new_n651_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n449_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n650_), .B1(new_n663_), .B2(new_n203_), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n478_), .A2(new_n479_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n486_), .A2(new_n204_), .A3(new_n666_), .A4(new_n646_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n661_), .A2(new_n583_), .A3(new_n666_), .A4(new_n651_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G8gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT108), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n668_), .A2(new_n672_), .A3(G8gat), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n670_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n671_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n667_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT40), .B(new_n667_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1325gat));
  INV_X1    g479(.A(G15gat), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n486_), .A2(new_n681_), .A3(new_n453_), .A4(new_n646_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n652_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT41), .B1(new_n684_), .B2(G15gat), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n683_), .A2(new_n686_), .A3(new_n681_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n682_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT109), .B(new_n682_), .C1(new_n685_), .C2(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1326gat));
  AOI21_X1  g491(.A(new_n394_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n693_));
  INV_X1    g492(.A(G22gat), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT42), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT42), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n482_), .A2(new_n694_), .ZN(new_n698_));
  OAI22_X1  g497(.A1(new_n696_), .A2(new_n697_), .B1(new_n647_), .B2(new_n698_), .ZN(G1327gat));
  NOR2_X1   g498(.A1(new_n583_), .A2(new_n610_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n645_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n486_), .A2(KEYINPUT112), .A3(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n238_), .B(new_n702_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT112), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n703_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G29gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n448_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n587_), .B(new_n710_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n588_), .B1(new_n476_), .B2(new_n485_), .ZN(new_n712_));
  XOR2_X1   g511(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n644_), .A2(new_n609_), .A3(new_n238_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n714_), .A2(KEYINPUT44), .A3(new_n716_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n448_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n721_), .B2(G29gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n709_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  INV_X1    g525(.A(G36gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n587_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n713_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n718_), .B(new_n715_), .C1(new_n730_), .C2(new_n711_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT44), .B1(new_n714_), .B2(new_n716_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n727_), .B1(new_n733_), .B2(new_n666_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n703_), .A2(new_n706_), .A3(new_n727_), .A4(new_n666_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n726_), .B1(new_n734_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n719_), .A2(new_n720_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G36gat), .B1(new_n739_), .B2(new_n665_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n735_), .B(KEYINPUT45), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(KEYINPUT46), .A3(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(G1329gat));
  INV_X1    g542(.A(G43gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n652_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n733_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n703_), .A2(new_n706_), .A3(new_n453_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n744_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n748_), .A3(new_n744_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n746_), .B(new_n747_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n750_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n719_), .A2(new_n720_), .A3(new_n745_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT47), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1330gat));
  OAI21_X1  g555(.A(G50gat), .B1(new_n739_), .B2(new_n394_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n394_), .A2(G50gat), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT114), .Z(new_n759_));
  NAND2_X1  g558(.A1(new_n707_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(G1331gat));
  AOI21_X1  g560(.A(new_n238_), .B1(new_n476_), .B2(new_n485_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n611_), .A2(new_n644_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G57gat), .B1(new_n765_), .B2(new_n448_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n661_), .A2(new_n583_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n609_), .A2(new_n238_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n645_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n449_), .A2(KEYINPUT115), .ZN(new_n771_));
  MUX2_X1   g570(.A(KEYINPUT115), .B(new_n771_), .S(G57gat), .Z(new_n772_));
  AOI21_X1  g571(.A(new_n766_), .B1(new_n770_), .B2(new_n772_), .ZN(G1332gat));
  INV_X1    g572(.A(new_n770_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G64gat), .B1(new_n774_), .B2(new_n665_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT48), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n665_), .A2(G64gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n764_), .B2(new_n777_), .ZN(G1333gat));
  OAI21_X1  g577(.A(G71gat), .B1(new_n774_), .B2(new_n652_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT49), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n652_), .A2(G71gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n764_), .B2(new_n781_), .ZN(G1334gat));
  OAI21_X1  g581(.A(G78gat), .B1(new_n774_), .B2(new_n394_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT50), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n394_), .A2(G78gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n764_), .B2(new_n785_), .ZN(G1335gat));
  NOR3_X1   g585(.A1(new_n644_), .A2(new_n610_), .A3(new_n238_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n714_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G85gat), .B1(new_n788_), .B2(new_n449_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n644_), .A2(new_n701_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n762_), .A2(new_n790_), .ZN(new_n791_));
  OR3_X1    g590(.A1(new_n791_), .A2(G85gat), .A3(new_n449_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n792_), .ZN(G1336gat));
  OAI21_X1  g592(.A(G92gat), .B1(new_n788_), .B2(new_n665_), .ZN(new_n794_));
  OR3_X1    g593(.A1(new_n791_), .A2(G92gat), .A3(new_n665_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n788_), .B2(new_n652_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n652_), .A2(new_n504_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n791_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(G1338gat));
  NAND4_X1  g600(.A1(new_n762_), .A2(new_n528_), .A3(new_n482_), .A4(new_n790_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n714_), .A2(new_n482_), .A3(new_n787_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n528_), .B1(new_n804_), .B2(KEYINPUT52), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(KEYINPUT52), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n803_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n802_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT53), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n802_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1339gat));
  NOR3_X1   g612(.A1(new_n652_), .A2(new_n395_), .A3(new_n449_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n816_));
  INV_X1    g615(.A(new_n583_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n540_), .A2(new_n613_), .ZN(new_n818_));
  AND4_X1   g617(.A1(new_n615_), .A2(new_n619_), .A3(new_n818_), .A4(new_n621_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n621_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n619_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n623_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n819_), .B1(new_n822_), .B2(KEYINPUT55), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n614_), .A2(KEYINPUT55), .A3(new_n615_), .A4(new_n619_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n628_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n615_), .B1(new_n614_), .B2(new_n619_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n620_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n629_), .B1(new_n831_), .B2(new_n824_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n828_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n238_), .A2(new_n630_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n827_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n223_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT120), .B(new_n218_), .C1(new_n220_), .C2(new_n222_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n225_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n237_), .B1(new_n232_), .B2(new_n224_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n233_), .A2(new_n237_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n817_), .B1(new_n837_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n826_), .A2(KEYINPUT56), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n843_), .A2(new_n630_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT121), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n843_), .A2(new_n630_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n832_), .A2(new_n828_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n848_), .A2(new_n853_), .A3(new_n854_), .A4(KEYINPUT58), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n587_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n831_), .A2(new_n824_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n828_), .B1(new_n857_), .B2(new_n628_), .ZN(new_n858_));
  AOI211_X1 g657(.A(KEYINPUT56), .B(new_n629_), .C1(new_n831_), .C2(new_n824_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT58), .B1(new_n860_), .B2(new_n853_), .ZN(new_n861_));
  OAI22_X1  g660(.A1(new_n847_), .A2(KEYINPUT57), .B1(new_n856_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863_));
  AOI211_X1 g662(.A(new_n863_), .B(new_n817_), .C1(new_n837_), .C2(new_n846_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n816_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n826_), .A2(KEYINPUT119), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n835_), .B1(new_n866_), .B2(new_n828_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n845_), .B1(new_n867_), .B2(new_n827_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n863_), .B1(new_n868_), .B2(new_n817_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n847_), .A2(KEYINPUT57), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n848_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n587_), .A3(new_n855_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n869_), .A2(KEYINPUT122), .A3(new_n870_), .A4(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n865_), .A2(new_n609_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n643_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n768_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT118), .B1(new_n644_), .B2(new_n768_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n588_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT54), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n881_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n644_), .A2(KEYINPUT118), .A3(new_n768_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n588_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n885_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n815_), .B1(new_n876_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(G113gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(new_n238_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n892_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n609_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n889_), .B1(new_n888_), .B2(new_n588_), .ZN(new_n897_));
  AOI211_X1 g696(.A(KEYINPUT54), .B(new_n587_), .C1(new_n886_), .C2(new_n887_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n814_), .B2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n901_), .B2(new_n814_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n895_), .A2(KEYINPUT59), .B1(new_n899_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n238_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n894_), .B1(new_n906_), .B2(new_n893_), .ZN(G1340gat));
  NAND2_X1  g706(.A1(new_n899_), .A2(new_n903_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n645_), .B(new_n908_), .C1(new_n892_), .C2(new_n900_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G120gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n644_), .A2(KEYINPUT60), .ZN(new_n911_));
  MUX2_X1   g710(.A(new_n911_), .B(KEYINPUT60), .S(G120gat), .Z(new_n912_));
  NAND2_X1  g711(.A1(new_n892_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n910_), .A2(KEYINPUT124), .A3(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1341gat));
  INV_X1    g717(.A(G127gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n892_), .A2(new_n919_), .A3(new_n610_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n904_), .A2(new_n610_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n922_), .B2(new_n919_), .ZN(G1342gat));
  INV_X1    g722(.A(G134gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n892_), .A2(new_n924_), .A3(new_n817_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n904_), .A2(new_n587_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n925_), .B1(new_n927_), .B2(new_n924_), .ZN(G1343gat));
  NAND2_X1  g727(.A1(new_n876_), .A2(new_n891_), .ZN(new_n929_));
  NOR4_X1   g728(.A1(new_n666_), .A2(new_n449_), .A3(new_n453_), .A4(new_n394_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n238_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n645_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g735(.A1(new_n931_), .A2(new_n609_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT61), .B(G155gat), .Z(new_n938_));
  XNOR2_X1  g737(.A(new_n937_), .B(new_n938_), .ZN(G1346gat));
  OR3_X1    g738(.A1(new_n931_), .A2(G162gat), .A3(new_n583_), .ZN(new_n940_));
  OAI21_X1  g739(.A(G162gat), .B1(new_n931_), .B2(new_n588_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1347gat));
  NOR3_X1   g741(.A1(new_n450_), .A2(new_n665_), .A3(new_n482_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n899_), .A2(new_n238_), .A3(new_n943_), .ZN(new_n944_));
  OAI21_X1  g743(.A(KEYINPUT62), .B1(new_n944_), .B2(KEYINPUT22), .ZN(new_n945_));
  OAI21_X1  g744(.A(G169gat), .B1(new_n944_), .B2(KEYINPUT62), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n947_), .B1(new_n279_), .B2(new_n945_), .ZN(G1348gat));
  AOI21_X1  g747(.A(new_n665_), .B1(new_n876_), .B2(new_n891_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n450_), .A2(new_n482_), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n949_), .A2(G176gat), .A3(new_n645_), .A4(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n951_), .A2(new_n952_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n899_), .A2(new_n943_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n955_), .A2(new_n644_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n956_), .A2(G176gat), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n953_), .A2(new_n954_), .A3(new_n957_), .ZN(G1349gat));
  NOR3_X1   g757(.A1(new_n955_), .A2(new_n260_), .A3(new_n609_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n949_), .A2(new_n610_), .A3(new_n950_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n960_), .A2(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n962_), .A2(G183gat), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n960_), .A2(new_n961_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n959_), .B1(new_n963_), .B2(new_n964_), .ZN(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n955_), .B2(new_n588_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n817_), .A2(new_n300_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n955_), .B2(new_n967_), .ZN(G1351gat));
  NOR2_X1   g767(.A1(new_n453_), .A2(new_n480_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n949_), .A2(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n971_), .A2(new_n238_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g772(.A1(new_n971_), .A2(new_n645_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g774(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n976_), .B1(new_n970_), .B2(new_n609_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n977_), .A2(KEYINPUT127), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979_));
  OAI211_X1 g778(.A(new_n979_), .B(new_n976_), .C1(new_n970_), .C2(new_n609_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n970_), .A2(new_n609_), .ZN(new_n981_));
  XOR2_X1   g780(.A(KEYINPUT63), .B(G211gat), .Z(new_n982_));
  AOI22_X1  g781(.A1(new_n978_), .A2(new_n980_), .B1(new_n981_), .B2(new_n982_), .ZN(G1354gat));
  OAI21_X1  g782(.A(G218gat), .B1(new_n970_), .B2(new_n588_), .ZN(new_n984_));
  OR2_X1    g783(.A1(new_n583_), .A2(G218gat), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n984_), .B1(new_n970_), .B2(new_n985_), .ZN(G1355gat));
endmodule


