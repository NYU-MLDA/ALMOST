//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202_));
  NAND3_X1  g001(.A1(new_n202_), .A2(G183gat), .A3(G190gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT83), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT23), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(G169gat), .B2(G176gat), .ZN(new_n210_));
  NOR3_X1   g009(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n213_), .A2(KEYINPUT82), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(KEYINPUT82), .ZN(new_n215_));
  OAI21_X1  g014(.A(G190gat), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n206_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n213_), .B2(G190gat), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n208_), .A2(new_n212_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n207_), .A2(new_n203_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(G183gat), .B2(G190gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(G169gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT30), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(G15gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(G71gat), .ZN(new_n234_));
  INV_X1    g033(.A(G99gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n230_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT87), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n237_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT85), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n242_), .B(new_n243_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(new_n245_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT84), .B(G43gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n241_), .B(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G225gat), .A2(G233gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT2), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT3), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  AOI211_X1 g068(.A(new_n258_), .B(new_n269_), .C1(KEYINPUT1), .C2(new_n265_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n248_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n268_), .A2(new_n273_), .A3(new_n247_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(KEYINPUT96), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT96), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n248_), .A2(new_n278_), .A3(new_n274_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n255_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n275_), .A2(KEYINPUT4), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n254_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n253_), .A3(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G29gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G85gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G57gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n282_), .A2(new_n290_), .A3(new_n283_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(KEYINPUT102), .A3(new_n291_), .ZN(new_n292_));
  AOI211_X1 g091(.A(KEYINPUT102), .B(new_n290_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n252_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G226gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT19), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT89), .B(G197gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT90), .B(G204gat), .ZN(new_n300_));
  OAI22_X1  g099(.A1(new_n299_), .A2(G204gat), .B1(new_n300_), .B2(G197gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT21), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(G204gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT21), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(G197gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G211gat), .B(G218gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n305_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n307_), .A2(new_n304_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT20), .B1(new_n312_), .B2(new_n228_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n226_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n217_), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT26), .B(G190gat), .Z(new_n317_));
  OAI211_X1 g116(.A(new_n212_), .B(new_n223_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n315_), .A2(new_n318_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n298_), .B1(new_n313_), .B2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G8gat), .B(G36gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT93), .ZN(new_n322_));
  XOR2_X1   g121(.A(G64gat), .B(G92gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT94), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n322_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n315_), .A2(new_n308_), .A3(new_n311_), .A4(new_n318_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n312_), .A2(new_n228_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n298_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT20), .A4(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n320_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT103), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n333_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n313_), .A2(new_n319_), .A3(new_n298_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n328_), .A2(KEYINPUT20), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT101), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n328_), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n329_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n341_), .B2(new_n298_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n334_), .B(new_n335_), .C1(new_n342_), .C2(new_n327_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT27), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT95), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n332_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n320_), .A2(new_n331_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n327_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n320_), .A2(new_n327_), .A3(KEYINPUT95), .A4(new_n331_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(KEYINPUT27), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n274_), .A2(KEYINPUT29), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n355_), .B(KEYINPUT28), .Z(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT91), .A2(G228gat), .A3(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G106gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n274_), .A2(KEYINPUT29), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n312_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G78gat), .ZN(new_n363_));
  AND2_X1   g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n364_), .A2(KEYINPUT91), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n360_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(new_n365_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G78gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n366_), .A3(G106gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G22gat), .B(G50gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n369_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n359_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n358_), .A3(new_n375_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n354_), .A2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n296_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n327_), .A2(KEYINPUT32), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n342_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n320_), .A3(new_n331_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n385_), .A2(new_n292_), .A3(new_n294_), .A4(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n289_), .A2(KEYINPUT98), .A3(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n346_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT98), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n290_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(KEYINPUT33), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n277_), .A2(new_n279_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n253_), .B1(new_n394_), .B2(KEYINPUT99), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(KEYINPUT99), .B2(new_n394_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n280_), .A2(new_n281_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT100), .B1(new_n397_), .B2(new_n253_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT100), .ZN(new_n399_));
  NOR4_X1   g198(.A1(new_n280_), .A2(new_n399_), .A3(new_n254_), .A4(new_n281_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n290_), .B(new_n396_), .C1(new_n398_), .C2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n389_), .A2(new_n390_), .A3(new_n393_), .A4(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n392_), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT97), .B1(new_n392_), .B2(KEYINPUT33), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n387_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n381_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n295_), .A2(new_n380_), .A3(new_n378_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n352_), .B1(KEYINPUT27), .B2(new_n343_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT104), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n378_), .A2(new_n380_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT104), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n354_), .A2(new_n411_), .A3(new_n412_), .A4(new_n295_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n407_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n252_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n383_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G29gat), .B(G36gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G43gat), .B(G50gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT80), .ZN(new_n420_));
  INV_X1    g219(.A(G1gat), .ZN(new_n421_));
  INV_X1    g220(.A(G8gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT14), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT77), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n424_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G15gat), .B(G22gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G8gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n425_), .A2(new_n431_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n420_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n419_), .B(KEYINPUT15), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n433_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G229gat), .A2(G233gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n420_), .B(new_n433_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G113gat), .B(G141gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G169gat), .B(G197gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  XNOR2_X1  g244(.A(new_n442_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT79), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n433_), .A2(G231gat), .A3(G233gat), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n433_), .B1(G231gat), .B2(G233gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G57gat), .B(G64gat), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(KEYINPUT11), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(KEYINPUT11), .ZN(new_n453_));
  XOR2_X1   g252(.A(G71gat), .B(G78gat), .Z(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n453_), .A2(new_n454_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OR3_X1    g256(.A1(new_n449_), .A2(new_n450_), .A3(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n457_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT78), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G127gat), .B(G155gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT16), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G183gat), .B(G211gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n458_), .A2(new_n459_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(KEYINPUT17), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n466_), .A2(KEYINPUT17), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n462_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n462_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n448_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n469_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n461_), .A3(new_n460_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n462_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(KEYINPUT79), .A3(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G190gat), .B(G218gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT75), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G134gat), .B(G162gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(KEYINPUT36), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT10), .B(G99gat), .ZN(new_n483_));
  OR3_X1    g282(.A1(new_n483_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT64), .B1(new_n483_), .B2(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G85gat), .ZN(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT9), .A3(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(KEYINPUT9), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT6), .B1(new_n235_), .B2(new_n360_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(G99gat), .A3(G106gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n486_), .A2(new_n491_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT7), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n499_), .B(new_n500_), .C1(G99gat), .C2(G106gat), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n235_), .B(new_n360_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n493_), .A2(new_n495_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT67), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n489_), .A2(new_n490_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n489_), .A2(KEYINPUT66), .A3(new_n490_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n498_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n512_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n501_), .A2(new_n502_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n515_), .A2(new_n516_), .A3(KEYINPUT8), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n497_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n435_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n503_), .A2(new_n504_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n515_), .B1(new_n520_), .B2(new_n507_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n513_), .A2(new_n498_), .ZN(new_n522_));
  OAI22_X1  g321(.A1(new_n521_), .A2(new_n498_), .B1(new_n522_), .B2(new_n516_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(new_n419_), .A3(new_n497_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G232gat), .A2(G233gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(KEYINPUT34), .Z(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  NAND3_X1  g327(.A1(new_n519_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n519_), .A2(new_n524_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n526_), .A2(new_n527_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n482_), .B(new_n529_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT76), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n532_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT74), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n541_), .A2(KEYINPUT76), .A3(new_n482_), .A4(new_n529_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n529_), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n481_), .B(KEYINPUT36), .Z(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(KEYINPUT37), .A3(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n477_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT70), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n457_), .B(new_n497_), .C1(new_n514_), .C2(new_n517_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G230gat), .A2(G233gat), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n555_), .A2(KEYINPUT69), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT69), .B1(new_n555_), .B2(new_n556_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n457_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT12), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n508_), .A2(new_n513_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n517_), .B1(new_n564_), .B2(KEYINPUT8), .ZN(new_n565_));
  INV_X1    g364(.A(new_n497_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n560_), .B(new_n563_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n457_), .B1(new_n523_), .B2(new_n497_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n554_), .B1(new_n559_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n556_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n555_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n572_), .B1(new_n568_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n555_), .A2(new_n556_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT69), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n555_), .A2(KEYINPUT69), .A3(new_n556_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n518_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n569_), .B1(new_n518_), .B2(new_n560_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n582_), .A3(KEYINPUT70), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n571_), .A2(new_n574_), .A3(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT72), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G120gat), .B(G148gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n584_), .A2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n571_), .A2(new_n583_), .A3(new_n574_), .A4(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT13), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR4_X1   g395(.A1(new_n416_), .A2(new_n447_), .A3(new_n553_), .A4(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n295_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n421_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n600_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n414_), .A2(new_n415_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n383_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n547_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n470_), .A2(new_n471_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n595_), .A2(new_n446_), .A3(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n421_), .B1(new_n609_), .B2(new_n598_), .ZN(new_n610_));
  OR3_X1    g409(.A1(new_n601_), .A2(new_n602_), .A3(new_n610_), .ZN(G1324gat));
  NAND3_X1  g410(.A1(new_n597_), .A2(new_n422_), .A3(new_n409_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n409_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n614_), .B2(G8gat), .ZN(new_n615_));
  AOI211_X1 g414(.A(KEYINPUT39), .B(new_n422_), .C1(new_n609_), .C2(new_n409_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(KEYINPUT40), .B(new_n612_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1325gat));
  AOI21_X1  g420(.A(new_n232_), .B1(new_n609_), .B2(new_n252_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT41), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n597_), .A2(new_n232_), .A3(new_n252_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n597_), .A2(new_n626_), .A3(new_n411_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n609_), .B2(new_n411_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(G1327gat));
  NOR2_X1   g431(.A1(new_n416_), .A2(new_n447_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n547_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n477_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(new_n596_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(G29gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n598_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n605_), .A2(new_n551_), .A3(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n543_), .A2(KEYINPUT37), .A3(new_n546_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT37), .B1(new_n543_), .B2(new_n546_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n640_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n646_));
  OAI22_X1  g445(.A1(new_n416_), .A2(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n641_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n595_), .A2(new_n477_), .A3(new_n446_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT44), .B1(new_n648_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n654_), .B(new_n651_), .C1(new_n641_), .C2(new_n647_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  AOI211_X1 g455(.A(KEYINPUT108), .B(new_n638_), .C1(new_n656_), .C2(new_n598_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n658_));
  INV_X1    g457(.A(new_n653_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n652_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n598_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n658_), .B1(new_n661_), .B2(G29gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n639_), .B1(new_n657_), .B2(new_n662_), .ZN(G1328gat));
  INV_X1    g462(.A(KEYINPUT46), .ZN(new_n664_));
  INV_X1    g463(.A(G36gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n656_), .B2(new_n409_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n354_), .A2(G36gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n633_), .A2(new_n636_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT109), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT109), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n633_), .A2(new_n670_), .A3(new_n636_), .A4(new_n667_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT45), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(KEYINPUT45), .A3(new_n671_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n664_), .B1(new_n666_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n674_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n672_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n653_), .A2(new_n655_), .A3(new_n354_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n678_), .B(KEYINPUT46), .C1(new_n679_), .C2(new_n665_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(G1329gat));
  AND2_X1   g480(.A1(new_n252_), .A2(G43gat), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n659_), .A2(new_n660_), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G43gat), .B1(new_n637_), .B2(new_n252_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT47), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n656_), .B2(new_n682_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(G1330gat));
  AND2_X1   g488(.A1(new_n411_), .A2(G50gat), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n659_), .A2(new_n660_), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G50gat), .B1(new_n637_), .B2(new_n411_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT110), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n656_), .B2(new_n690_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1331gat));
  NAND2_X1  g496(.A1(new_n472_), .A2(new_n476_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n595_), .A2(new_n446_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n605_), .A2(new_n547_), .A3(new_n698_), .A4(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G57gat), .B1(new_n700_), .B2(new_n295_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n552_), .A2(new_n596_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT111), .Z(new_n703_));
  NOR2_X1   g502(.A1(new_n416_), .A2(new_n446_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n295_), .A2(G57gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n701_), .B1(new_n705_), .B2(new_n706_), .ZN(G1332gat));
  INV_X1    g506(.A(G64gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n700_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n409_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n710_), .A2(new_n711_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n409_), .A2(new_n708_), .ZN(new_n714_));
  OAI22_X1  g513(.A1(new_n712_), .A2(new_n713_), .B1(new_n705_), .B2(new_n714_), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n700_), .B2(new_n415_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT49), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n415_), .A2(G71gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n705_), .B2(new_n718_), .ZN(G1334gat));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n709_), .A2(new_n411_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G78gat), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT50), .B(new_n363_), .C1(new_n709_), .C2(new_n411_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n411_), .A2(new_n363_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT113), .Z(new_n725_));
  OAI22_X1  g524(.A1(new_n722_), .A2(new_n723_), .B1(new_n705_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT114), .ZN(G1335gat));
  NOR4_X1   g526(.A1(new_n416_), .A2(new_n446_), .A3(new_n595_), .A4(new_n635_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(new_n487_), .A3(new_n598_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n699_), .A2(new_n477_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n645_), .A2(new_n646_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n605_), .B2(new_n551_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n416_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT115), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n648_), .A2(KEYINPUT115), .A3(new_n731_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n295_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n729_), .B1(new_n739_), .B2(new_n487_), .ZN(G1336gat));
  AOI21_X1  g539(.A(G92gat), .B1(new_n728_), .B2(new_n409_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT116), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n737_), .A2(new_n738_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n354_), .A2(new_n488_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n743_), .B2(new_n744_), .ZN(G1337gat));
  INV_X1    g544(.A(new_n483_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n728_), .A2(new_n252_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n415_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n235_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT51), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n747_), .C1(new_n748_), .C2(new_n235_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n728_), .A2(new_n360_), .A3(new_n411_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n648_), .A2(new_n411_), .A3(new_n731_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(G106gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G106gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n754_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  INV_X1    g562(.A(G113gat), .ZN(new_n764_));
  INV_X1    g563(.A(new_n607_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n441_), .A2(new_n439_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n766_), .B(new_n445_), .C1(new_n439_), .C2(new_n437_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n437_), .A2(KEYINPUT118), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n768_), .A2(new_n438_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n445_), .B1(new_n441_), .B2(new_n438_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n767_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(new_n593_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n571_), .A2(new_n777_), .A3(new_n583_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n570_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n567_), .B(new_n555_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n779_), .A2(KEYINPUT55), .B1(new_n572_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n782_), .B2(new_n591_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n784_), .B(new_n590_), .C1(new_n778_), .C2(new_n781_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n776_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT58), .B(new_n776_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n551_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n594_), .B2(new_n775_), .ZN(new_n792_));
  AOI211_X1 g591(.A(KEYINPUT119), .B(new_n774_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n446_), .B(new_n593_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n634_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n790_), .B1(new_n796_), .B2(KEYINPUT57), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n798_), .B(new_n634_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n765_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n552_), .A2(new_n447_), .A3(new_n595_), .A4(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n644_), .A2(new_n595_), .A3(new_n447_), .A4(new_n698_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n801_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n800_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n382_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n415_), .A2(new_n295_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n594_), .A2(new_n775_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT119), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n594_), .A2(new_n791_), .A3(new_n775_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n446_), .A2(new_n593_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n782_), .A2(new_n591_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n784_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n782_), .A2(KEYINPUT56), .A3(new_n591_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n815_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n547_), .B1(new_n814_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n798_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n796_), .A2(KEYINPUT57), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n790_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n477_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n806_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n809_), .A2(new_n808_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(KEYINPUT59), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n810_), .A2(KEYINPUT59), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n764_), .B1(new_n828_), .B2(new_n446_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n810_), .A2(G113gat), .A3(new_n447_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT120), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(new_n827_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n802_), .A2(new_n805_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n823_), .B2(new_n765_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n826_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837_), .B2(new_n447_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  INV_X1    g638(.A(new_n830_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n831_), .A2(new_n841_), .ZN(G1340gat));
  XOR2_X1   g641(.A(KEYINPUT121), .B(G120gat), .Z(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n595_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n835_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n843_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n837_), .A2(new_n595_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n843_), .ZN(G1341gat));
  AOI21_X1  g646(.A(G127gat), .B1(new_n835_), .B2(new_n698_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT122), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n607_), .A2(G127gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n828_), .B2(new_n850_), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n828_), .B2(new_n551_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n810_), .A2(G134gat), .A3(new_n547_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT123), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G134gat), .B1(new_n837_), .B2(new_n644_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857_));
  INV_X1    g656(.A(new_n854_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n859_), .ZN(G1343gat));
  NAND4_X1  g659(.A1(new_n415_), .A2(new_n354_), .A3(new_n411_), .A4(new_n598_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT124), .B1(new_n834_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n863_));
  INV_X1    g662(.A(new_n861_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n551_), .A2(new_n789_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n820_), .A2(new_n798_), .B1(new_n865_), .B2(new_n788_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n607_), .B1(new_n866_), .B2(new_n822_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n863_), .B(new_n864_), .C1(new_n867_), .C2(new_n833_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n862_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n446_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n596_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT125), .B(G148gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1345gat));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n869_), .B2(new_n698_), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n477_), .B(new_n875_), .C1(new_n862_), .C2(new_n868_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n877_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n863_), .B1(new_n807_), .B2(new_n864_), .ZN(new_n882_));
  AOI211_X1 g681(.A(KEYINPUT124), .B(new_n861_), .C1(new_n800_), .C2(new_n806_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n698_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n875_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n869_), .A2(new_n698_), .A3(new_n876_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n879_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n881_), .A2(new_n887_), .ZN(G1346gat));
  INV_X1    g687(.A(new_n869_), .ZN(new_n889_));
  OR3_X1    g688(.A1(new_n889_), .A2(G162gat), .A3(new_n547_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G162gat), .B1(new_n889_), .B2(new_n644_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1347gat));
  NOR3_X1   g691(.A1(new_n296_), .A2(new_n354_), .A3(new_n411_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n825_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n446_), .ZN(new_n895_));
  OAI211_X1 g694(.A(KEYINPUT62), .B(G169gat), .C1(new_n895_), .C2(KEYINPUT22), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  INV_X1    g696(.A(new_n895_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT22), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(G169gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n898_), .B2(new_n897_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n896_), .B1(new_n900_), .B2(new_n902_), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n894_), .B2(new_n596_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n807_), .A2(new_n893_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n596_), .A2(G176gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1349gat));
  AOI21_X1  g706(.A(G183gat), .B1(new_n905_), .B2(new_n698_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n765_), .A2(new_n217_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n894_), .B2(new_n909_), .ZN(G1350gat));
  NOR2_X1   g709(.A1(new_n547_), .A2(new_n317_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n894_), .A2(new_n911_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n894_), .A2(new_n551_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n206_), .ZN(G1351gat));
  NOR4_X1   g713(.A1(new_n834_), .A2(new_n354_), .A3(new_n252_), .A4(new_n408_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n446_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n596_), .ZN(new_n918_));
  MUX2_X1   g717(.A(new_n300_), .B(G204gat), .S(new_n918_), .Z(G1353gat));
  NAND2_X1  g718(.A1(new_n915_), .A2(new_n607_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  AND2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n920_), .B2(new_n921_), .ZN(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n915_), .A2(new_n925_), .A3(new_n634_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n915_), .A2(new_n551_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n925_), .ZN(G1355gat));
endmodule


