//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n978_, new_n979_, new_n981_, new_n982_, new_n984_, new_n985_,
    new_n986_, new_n988_, new_n989_, new_n990_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_;
  NAND3_X1  g000(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT87), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT87), .ZN(new_n204_));
  NAND4_X1  g003(.A1(new_n204_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207_));
  INV_X1    g006(.A(G141gat), .ZN(new_n208_));
  INV_X1    g007(.A(G148gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT88), .B1(new_n206_), .B2(new_n215_), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n203_), .A2(new_n205_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n223_), .A2(KEYINPUT86), .A3(KEYINPUT1), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT86), .B1(new_n223_), .B2(KEYINPUT1), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(KEYINPUT1), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n227_), .A2(new_n222_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n230_), .A2(new_n232_), .A3(new_n211_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n226_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT28), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT28), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n226_), .A2(new_n238_), .A3(new_n235_), .A4(new_n234_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G22gat), .B(G50gat), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G78gat), .B(G106gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT92), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n224_), .B1(new_n216_), .B2(new_n220_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT29), .B1(new_n247_), .B2(new_n233_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(KEYINPUT89), .B(KEYINPUT29), .C1(new_n247_), .C2(new_n233_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G211gat), .B(G218gat), .Z(new_n252_));
  OR2_X1    g051(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n253_));
  INV_X1    g052(.A(G204gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT21), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(G197gat), .B2(G204gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n252_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n254_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G197gat), .A2(G204gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(KEYINPUT21), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(KEYINPUT21), .A3(new_n252_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G228gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n250_), .A2(new_n251_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT91), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n263_), .A2(new_n264_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n248_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n269_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n270_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n246_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n248_), .A2(new_n271_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n267_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT91), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n279_), .A2(new_n245_), .A3(new_n274_), .A4(new_n269_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n243_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n274_), .A3(new_n269_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT93), .B1(new_n282_), .B2(new_n244_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n243_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(KEYINPUT93), .A3(new_n244_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n281_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT26), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(G190gat), .ZN(new_n289_));
  INV_X1    g088(.A(G190gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(KEYINPUT26), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT95), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G183gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT25), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G183gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(KEYINPUT26), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n288_), .A2(G190gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT95), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n292_), .A2(new_n297_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(G169gat), .B2(G176gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT96), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT96), .B1(new_n308_), .B2(new_n303_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n306_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT97), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n302_), .A2(new_n312_), .A3(KEYINPUT97), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT23), .B1(new_n293_), .B2(new_n290_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G183gat), .A3(G190gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(KEYINPUT83), .B(KEYINPUT23), .C1(new_n293_), .C2(new_n290_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n310_), .A2(new_n303_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n315_), .A2(new_n316_), .A3(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n317_), .A2(new_n319_), .A3(KEYINPUT81), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT81), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n328_), .A2(new_n318_), .A3(G183gat), .A4(G190gat), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n327_), .B(new_n329_), .C1(G183gat), .C2(G190gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT22), .B(G169gat), .ZN(new_n331_));
  INV_X1    g130(.A(G176gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n308_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n326_), .A2(new_n265_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n294_), .A2(new_n296_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n304_), .A2(new_n311_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n327_), .A2(new_n329_), .A3(new_n323_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(new_n338_), .A3(KEYINPUT80), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT82), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G169gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n345_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G169gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n321_), .A2(new_n322_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n347_), .B(new_n351_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n344_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n336_), .B1(new_n355_), .B2(new_n271_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n335_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT20), .B1(new_n355_), .B2(new_n271_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n302_), .A2(new_n312_), .A3(KEYINPUT97), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT97), .B1(new_n302_), .B2(new_n312_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n324_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n334_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n271_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n360_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n363_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n361_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G8gat), .B(G36gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT18), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n371_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n265_), .B1(new_n326_), .B2(new_n334_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n360_), .B1(new_n378_), .B2(new_n362_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n335_), .A2(new_n356_), .A3(new_n369_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n375_), .A3(new_n380_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n377_), .A2(KEYINPUT27), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n379_), .A2(new_n375_), .A3(new_n380_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n375_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT99), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n379_), .A2(new_n380_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n376_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n381_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(KEYINPUT99), .A3(new_n383_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n382_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G127gat), .B(G134gat), .Z(new_n394_));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT84), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G113gat), .B(G120gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n396_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n226_), .A2(new_n234_), .A3(new_n404_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n396_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n400_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n247_), .B2(new_n233_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n409_), .A3(KEYINPUT4), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n408_), .B(new_n411_), .C1(new_n247_), .C2(new_n233_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT98), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n405_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G85gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT0), .B(G57gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  NAND3_X1  g219(.A1(new_n415_), .A2(new_n416_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n287_), .B1(new_n393_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n408_), .B(KEYINPUT31), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G43gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n355_), .B(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(G15gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT30), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n429_), .B(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n426_), .B1(new_n435_), .B2(KEYINPUT85), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(KEYINPUT85), .B2(new_n435_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n435_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT85), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n426_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n282_), .A2(new_n244_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT93), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n280_), .A2(new_n243_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n286_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n281_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n375_), .A2(KEYINPUT32), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n371_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n379_), .A2(new_n380_), .A3(new_n449_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n451_), .B(new_n452_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n421_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n410_), .A2(new_n413_), .A3(new_n412_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n420_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n405_), .A2(new_n409_), .A3(new_n414_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n455_), .A2(new_n381_), .A3(new_n390_), .A4(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n421_), .A2(new_n454_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n453_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n441_), .B1(new_n448_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT100), .B1(new_n425_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n377_), .A2(KEYINPUT27), .A3(new_n381_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT99), .B1(new_n391_), .B2(new_n383_), .ZN(new_n466_));
  AOI211_X1 g265(.A(new_n387_), .B(KEYINPUT27), .C1(new_n390_), .C2(new_n381_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n424_), .B(new_n465_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n448_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT100), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n460_), .A2(new_n461_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n287_), .A2(new_n471_), .A3(new_n453_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n469_), .A2(new_n470_), .A3(new_n472_), .A4(new_n441_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n465_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT101), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT101), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n393_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n448_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n424_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n441_), .A2(new_n479_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n464_), .A2(new_n473_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(G22gat), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(G22gat), .B1(new_n486_), .B2(new_n487_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n485_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G1gat), .B(G8gat), .Z(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT73), .B(G15gat), .ZN(new_n495_));
  INV_X1    g294(.A(G22gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n488_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n492_), .A3(new_n485_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G29gat), .B(G36gat), .Z(new_n500_));
  XOR2_X1   g299(.A(G43gat), .B(G50gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G29gat), .B(G36gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n494_), .A2(new_n499_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n502_), .A2(KEYINPUT15), .A3(new_n505_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT15), .B1(new_n502_), .B2(new_n505_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n494_), .A2(new_n499_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT77), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n507_), .B(new_n508_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT76), .ZN(new_n517_));
  INV_X1    g316(.A(new_n506_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n498_), .A2(new_n492_), .A3(new_n485_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n492_), .B1(new_n498_), .B2(new_n485_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n507_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n508_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n517_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AOI211_X1 g323(.A(KEYINPUT76), .B(new_n508_), .C1(new_n521_), .C2(new_n507_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n516_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n482_), .B1(new_n526_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n526_), .A2(new_n482_), .A3(new_n530_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n516_), .B(new_n529_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT79), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n524_), .A2(new_n525_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT79), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n516_), .A4(new_n529_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n532_), .A2(new_n533_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G230gat), .A2(G233gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT10), .B(G99gat), .ZN(new_n543_));
  OR3_X1    g342(.A1(new_n543_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(G85gat), .B(G92gat), .Z(new_n545_));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT6), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(G99gat), .A3(G106gat), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n545_), .A2(KEYINPUT9), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT65), .B(G92gat), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(G85gat), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT64), .B1(new_n543_), .B2(G106gat), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n544_), .A2(new_n550_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT8), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(new_n549_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT67), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n559_));
  INV_X1    g358(.A(G99gat), .ZN(new_n560_));
  INV_X1    g359(.A(G106gat), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT67), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n547_), .A2(new_n549_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n558_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n556_), .B1(new_n568_), .B2(new_n545_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n556_), .A2(KEYINPUT66), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n556_), .A2(KEYINPUT66), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n545_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n557_), .B2(new_n565_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n555_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT11), .ZN(new_n576_));
  INV_X1    g375(.A(G57gat), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(G64gat), .ZN(new_n578_));
  INV_X1    g377(.A(G64gat), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(G57gat), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n576_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(G57gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(G64gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT11), .ZN(new_n584_));
  XOR2_X1   g383(.A(G71gat), .B(G78gat), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G71gat), .B(G78gat), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n587_), .A2(KEYINPUT11), .A3(new_n582_), .A4(new_n583_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n575_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n575_), .A3(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n574_), .A2(new_n592_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n586_), .A2(new_n575_), .A3(new_n588_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(new_n589_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n565_), .A2(new_n557_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n596_), .A2(new_n545_), .A3(new_n570_), .A4(new_n571_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n545_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n566_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n564_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n600_), .B2(new_n567_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n601_), .B2(new_n556_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n595_), .A2(new_n602_), .A3(new_n555_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n593_), .A2(new_n603_), .A3(KEYINPUT12), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT12), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n574_), .A2(new_n592_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n542_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n593_), .A2(new_n603_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n542_), .B2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(G120gat), .B(G148gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n604_), .A2(new_n606_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n541_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n542_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n614_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n540_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n609_), .A2(new_n615_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n614_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(KEYINPUT13), .A3(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n574_), .A2(new_n511_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT34), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n633_));
  OAI221_X1 g432(.A(new_n630_), .B1(new_n518_), .B2(new_n574_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(KEYINPUT36), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n639_), .B(KEYINPUT36), .Z(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n636_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n629_), .B1(new_n642_), .B2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n641_), .B(new_n628_), .C1(new_n636_), .C2(new_n644_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(G231gat), .ZN(new_n649_));
  INV_X1    g448(.A(G233gat), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n494_), .A2(new_n499_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n592_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n655_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n595_), .A3(new_n653_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT74), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(G127gat), .B(G155gat), .Z(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT16), .ZN(new_n662_));
  XNOR2_X1  g461(.A(G183gat), .B(G211gat), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n660_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n656_), .A2(new_n658_), .A3(new_n664_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT17), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT17), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n669_), .B(KEYINPUT75), .C1(new_n670_), .C2(new_n666_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT75), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n666_), .A2(new_n670_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(KEYINPUT17), .A2(new_n667_), .B1(new_n660_), .B2(new_n665_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n648_), .A2(new_n676_), .ZN(new_n677_));
  NOR4_X1   g476(.A1(new_n481_), .A2(new_n539_), .A3(new_n627_), .A4(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n678_), .A2(new_n483_), .A3(new_n479_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT38), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n539_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n626_), .A2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT102), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n673_), .A2(new_n674_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n642_), .A2(new_n645_), .ZN(new_n686_));
  NOR4_X1   g485(.A1(new_n481_), .A2(new_n684_), .A3(new_n685_), .A4(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n483_), .B1(new_n687_), .B2(new_n479_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n681_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n680_), .B2(new_n679_), .ZN(G1324gat));
  AND2_X1   g489(.A1(new_n475_), .A2(new_n477_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n678_), .A2(new_n484_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n687_), .A2(new_n691_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G8gat), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT39), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(KEYINPUT39), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1325gat));
  INV_X1    g498(.A(new_n441_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n431_), .B1(new_n687_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT41), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n678_), .A2(new_n431_), .A3(new_n700_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1326gat));
  NAND3_X1  g503(.A1(new_n678_), .A2(new_n496_), .A3(new_n448_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n687_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G22gat), .B1(new_n706_), .B2(new_n287_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT42), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT42), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT103), .ZN(G1327gat));
  NOR2_X1   g510(.A1(new_n481_), .A2(new_n539_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n676_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n686_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n627_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n716_), .A2(G29gat), .A3(new_n424_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n464_), .A2(new_n473_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n478_), .A2(new_n480_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n721_));
  INV_X1    g520(.A(new_n648_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n481_), .B2(new_n648_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n683_), .B(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n713_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT44), .B1(new_n725_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731_));
  AOI211_X1 g530(.A(new_n731_), .B(new_n728_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT104), .B1(new_n733_), .B2(new_n479_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n721_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n481_), .A2(KEYINPUT43), .A3(new_n648_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n729_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n731_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n725_), .A2(KEYINPUT44), .A3(new_n729_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n738_), .A2(KEYINPUT104), .A3(new_n479_), .A4(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G29gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n717_), .B1(new_n734_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT105), .B(new_n717_), .C1(new_n734_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1328gat));
  NAND2_X1  g545(.A1(new_n733_), .A2(new_n691_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G36gat), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(G36gat), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n691_), .A2(KEYINPUT106), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n691_), .A2(KEYINPUT106), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n712_), .A2(new_n753_), .A3(new_n715_), .A4(new_n756_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(KEYINPUT45), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT45), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n758_), .A2(new_n759_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n748_), .A2(new_n752_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n752_), .B1(new_n748_), .B2(new_n760_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1329gat));
  NAND3_X1  g562(.A1(new_n712_), .A2(new_n700_), .A3(new_n715_), .ZN(new_n764_));
  INV_X1    g563(.A(G43gat), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT109), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n441_), .A2(new_n765_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n738_), .A2(new_n739_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n738_), .A2(KEYINPUT108), .A3(new_n739_), .A4(new_n768_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n767_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n774_), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n776_), .B(new_n767_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1330gat));
  NAND3_X1  g577(.A1(new_n733_), .A2(G50gat), .A3(new_n448_), .ZN(new_n779_));
  INV_X1    g578(.A(G50gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n716_), .B2(new_n287_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1331gat));
  NOR4_X1   g581(.A1(new_n481_), .A2(new_n682_), .A3(new_n626_), .A4(new_n677_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n577_), .A3(new_n479_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n686_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n682_), .A2(new_n713_), .ZN(new_n786_));
  AND4_X1   g585(.A1(new_n720_), .A2(new_n627_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n479_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n788_), .B2(new_n577_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT111), .ZN(G1332gat));
  AOI21_X1  g589(.A(new_n579_), .B1(new_n787_), .B2(new_n756_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT48), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n783_), .A2(new_n579_), .A3(new_n756_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1333gat));
  INV_X1    g593(.A(G71gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n787_), .B2(new_n700_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT49), .Z(new_n797_));
  NAND3_X1  g596(.A1(new_n783_), .A2(new_n795_), .A3(new_n700_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1334gat));
  INV_X1    g598(.A(G78gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n787_), .B2(new_n448_), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT50), .Z(new_n802_));
  NAND3_X1  g601(.A1(new_n783_), .A2(new_n800_), .A3(new_n448_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1335gat));
  NOR4_X1   g603(.A1(new_n481_), .A2(new_n682_), .A3(new_n626_), .A4(new_n714_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT112), .ZN(new_n806_));
  AOI21_X1  g605(.A(G85gat), .B1(new_n806_), .B2(new_n479_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n626_), .A2(new_n682_), .A3(new_n676_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n725_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n479_), .A2(G85gat), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT113), .Z(new_n811_));
  AOI21_X1  g610(.A(new_n807_), .B1(new_n809_), .B2(new_n811_), .ZN(G1336gat));
  AOI21_X1  g611(.A(G92gat), .B1(new_n806_), .B2(new_n691_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n756_), .A2(new_n551_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n809_), .B2(new_n814_), .ZN(G1337gat));
  NOR2_X1   g614(.A1(new_n441_), .A2(new_n543_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n806_), .A2(new_n816_), .B1(new_n817_), .B2(KEYINPUT51), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n809_), .A2(new_n700_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G99gat), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n817_), .A2(KEYINPUT51), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n821_), .B(new_n822_), .Z(G1338gat));
  NAND3_X1  g622(.A1(new_n806_), .A2(new_n561_), .A3(new_n448_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n809_), .A2(new_n448_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(G106gat), .ZN(new_n827_));
  AOI211_X1 g626(.A(KEYINPUT52), .B(new_n561_), .C1(new_n809_), .C2(new_n448_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n824_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT53), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n824_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1339gat));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n478_), .A2(new_n479_), .A3(new_n700_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n533_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n531_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n538_), .A2(new_n535_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n623_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n618_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT116), .B1(new_n607_), .B2(KEYINPUT55), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n607_), .A2(KEYINPUT55), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n604_), .A2(new_n542_), .A3(new_n606_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .A4(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n614_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT56), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(KEYINPUT56), .A3(new_n614_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n841_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n538_), .A2(new_n535_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n529_), .B1(new_n522_), .B2(new_n508_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n514_), .A2(new_n515_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n507_), .A2(new_n523_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n854_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n623_), .A2(new_n624_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n785_), .B1(new_n853_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n623_), .A2(new_n854_), .A3(new_n858_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n848_), .A2(KEYINPUT56), .A3(new_n614_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT56), .B1(new_n848_), .B2(new_n614_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n648_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT58), .B(new_n866_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n864_), .A2(new_n863_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n865_), .B1(new_n873_), .B2(KEYINPUT117), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n863_), .A2(new_n864_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n872_), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n875_), .A2(KEYINPUT117), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n713_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n622_), .A2(new_n676_), .A3(new_n539_), .A4(new_n625_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n648_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n786_), .A2(new_n626_), .A3(KEYINPUT115), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n881_), .A4(new_n648_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n884_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n837_), .B1(new_n878_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n875_), .A2(new_n876_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n863_), .A2(new_n864_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n685_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n889_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n836_), .B1(new_n894_), .B2(new_n835_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n834_), .B1(new_n890_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n873_), .A2(new_n865_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n888_), .B1(new_n897_), .B2(new_n685_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n835_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT59), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n891_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n873_), .A2(KEYINPUT117), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n865_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n888_), .B1(new_n904_), .B2(new_n713_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n900_), .B(KEYINPUT118), .C1(new_n905_), .C2(new_n837_), .ZN(new_n906_));
  INV_X1    g705(.A(G113gat), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n539_), .A2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n896_), .A2(new_n906_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n894_), .A2(new_n835_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n907_), .B1(new_n910_), .B2(new_n539_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n909_), .A2(KEYINPUT119), .A3(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1340gat));
  OAI21_X1  g715(.A(new_n900_), .B1(new_n905_), .B2(new_n837_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G120gat), .B1(new_n917_), .B2(new_n626_), .ZN(new_n918_));
  INV_X1    g717(.A(G120gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n919_), .B1(new_n626_), .B2(KEYINPUT60), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(KEYINPUT60), .B2(new_n919_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n918_), .B1(new_n910_), .B2(new_n921_), .ZN(G1341gat));
  XOR2_X1   g721(.A(KEYINPUT120), .B(G127gat), .Z(new_n923_));
  NOR2_X1   g722(.A1(new_n685_), .A2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n896_), .A2(new_n906_), .A3(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(G127gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n910_), .B2(new_n713_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT121), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n925_), .A2(new_n930_), .A3(new_n927_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1342gat));
  NAND3_X1  g731(.A1(new_n896_), .A2(new_n722_), .A3(new_n906_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G134gat), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n785_), .A2(G134gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n910_), .B2(new_n935_), .ZN(G1343gat));
  NAND2_X1  g735(.A1(new_n448_), .A2(new_n441_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n898_), .A2(new_n937_), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n938_), .A2(new_n479_), .A3(new_n754_), .A4(new_n755_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n539_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(new_n208_), .ZN(G1344gat));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n626_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n209_), .ZN(G1345gat));
  NOR2_X1   g742(.A1(new_n939_), .A2(new_n713_), .ZN(new_n944_));
  XOR2_X1   g743(.A(KEYINPUT61), .B(G155gat), .Z(new_n945_));
  XNOR2_X1  g744(.A(new_n944_), .B(new_n945_), .ZN(G1346gat));
  INV_X1    g745(.A(G162gat), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n939_), .A2(new_n947_), .A3(new_n648_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n939_), .B2(new_n785_), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n949_), .A2(KEYINPUT122), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(KEYINPUT122), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n948_), .B1(new_n950_), .B2(new_n951_), .ZN(G1347gat));
  AOI21_X1  g751(.A(new_n479_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(new_n700_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(KEYINPUT123), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n953_), .A2(new_n956_), .A3(new_n700_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n448_), .B1(new_n955_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n878_), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n958_), .B(new_n682_), .C1(new_n959_), .C2(new_n888_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(G169gat), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n960_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n963_), .A2(KEYINPUT62), .A3(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(KEYINPUT124), .B1(new_n960_), .B2(G169gat), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967_));
  INV_X1    g766(.A(new_n960_), .ZN(new_n968_));
  AOI22_X1  g767(.A1(new_n966_), .A2(new_n967_), .B1(new_n331_), .B2(new_n968_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n965_), .A2(new_n969_), .ZN(G1348gat));
  AND2_X1   g769(.A1(new_n955_), .A2(new_n957_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n894_), .A2(new_n287_), .ZN(new_n972_));
  NOR4_X1   g771(.A1(new_n971_), .A2(new_n972_), .A3(new_n332_), .A4(new_n626_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n958_), .B1(new_n959_), .B2(new_n888_), .ZN(new_n974_));
  INV_X1    g773(.A(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(new_n627_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n973_), .B1(new_n976_), .B2(new_n332_), .ZN(G1349gat));
  NOR3_X1   g776(.A1(new_n974_), .A2(new_n297_), .A3(new_n685_), .ZN(new_n978_));
  OR3_X1    g777(.A1(new_n971_), .A2(new_n713_), .A3(new_n972_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n293_), .B2(new_n979_), .ZN(G1350gat));
  OAI21_X1  g779(.A(G190gat), .B1(new_n974_), .B2(new_n648_), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n686_), .A2(new_n292_), .A3(new_n301_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n974_), .B2(new_n982_), .ZN(G1351gat));
  NAND2_X1  g782(.A1(new_n938_), .A2(new_n953_), .ZN(new_n984_));
  INV_X1    g783(.A(new_n984_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n985_), .A2(new_n682_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n986_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988_));
  OAI211_X1 g787(.A(new_n985_), .B(new_n627_), .C1(new_n988_), .C2(new_n254_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n988_), .A2(new_n254_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n989_), .B(new_n990_), .ZN(G1353gat));
  NOR3_X1   g790(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992_));
  AND2_X1   g791(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n993_));
  NOR4_X1   g792(.A1(new_n984_), .A2(new_n685_), .A3(new_n992_), .A4(new_n993_), .ZN(new_n994_));
  OAI21_X1  g793(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n995_));
  XNOR2_X1  g794(.A(new_n994_), .B(new_n995_), .ZN(G1354gat));
  INV_X1    g795(.A(G218gat), .ZN(new_n997_));
  NAND3_X1  g796(.A1(new_n985_), .A2(new_n997_), .A3(new_n686_), .ZN(new_n998_));
  NOR2_X1   g797(.A1(new_n984_), .A2(new_n648_), .ZN(new_n999_));
  OAI21_X1  g798(.A(new_n998_), .B1(new_n997_), .B2(new_n999_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n1000_), .A2(KEYINPUT127), .ZN(new_n1001_));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1002_));
  OAI211_X1 g801(.A(new_n998_), .B(new_n1002_), .C1(new_n997_), .C2(new_n999_), .ZN(new_n1003_));
  NAND2_X1  g802(.A1(new_n1001_), .A2(new_n1003_), .ZN(G1355gat));
endmodule


