//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT26), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(G190gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT26), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n202_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT25), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT25), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT78), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT79), .B1(new_n203_), .B2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(new_n208_), .B2(G183gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n207_), .A2(new_n212_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT24), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT23), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n216_), .A2(KEYINPUT80), .A3(new_n220_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(new_n225_), .A3(new_n226_), .A4(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT82), .B(G169gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT81), .ZN(new_n231_));
  AOI21_X1  g030(.A(G176gat), .B1(new_n231_), .B2(KEYINPUT22), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n230_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n225_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT83), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n233_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n229_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT30), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT84), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G15gat), .B(G43gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G71gat), .B(G99gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT84), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n244_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n255_), .A3(KEYINPUT86), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G127gat), .B(G134gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G120gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT85), .B(G113gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT31), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n251_), .A2(new_n255_), .A3(KEYINPUT86), .A4(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n268_), .B1(G155gat), .B2(G162gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n270_), .A2(KEYINPUT87), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT1), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(KEYINPUT88), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n270_), .A2(KEYINPUT87), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n268_), .A2(G155gat), .A3(G162gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n276_), .B1(new_n280_), .B2(new_n273_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n277_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT89), .ZN(new_n284_));
  XOR2_X1   g083(.A(G141gat), .B(G148gat), .Z(new_n285_));
  AND3_X1   g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT90), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n288_), .B1(new_n289_), .B2(KEYINPUT2), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT2), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n291_), .A2(KEYINPUT90), .A3(G141gat), .A4(G148gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G141gat), .ZN(new_n294_));
  INV_X1    g093(.A(G148gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(KEYINPUT3), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(G141gat), .B2(G148gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n289_), .A2(KEYINPUT2), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n293_), .A2(new_n299_), .A3(KEYINPUT91), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n278_), .A2(new_n279_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n296_), .A2(new_n298_), .B1(new_n289_), .B2(KEYINPUT2), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT91), .B1(new_n304_), .B2(new_n293_), .ZN(new_n305_));
  NOR4_X1   g104(.A1(new_n303_), .A2(new_n305_), .A3(KEYINPUT92), .A4(new_n273_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT92), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n301_), .A2(new_n302_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n293_), .A2(new_n300_), .A3(new_n299_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT91), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n273_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n307_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  OAI22_X1  g111(.A1(new_n286_), .A2(new_n287_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT93), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n283_), .A2(new_n285_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT89), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n311_), .A2(new_n302_), .A3(new_n301_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT92), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n308_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n323_), .A3(KEYINPUT93), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n315_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n267_), .B1(new_n325_), .B2(KEYINPUT29), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n315_), .A2(new_n324_), .A3(new_n327_), .A4(new_n266_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G228gat), .A2(G233gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n313_), .A2(KEYINPUT29), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT95), .B(G197gat), .ZN(new_n333_));
  OAI211_X1 g132(.A(KEYINPUT21), .B(new_n332_), .C1(new_n333_), .C2(G204gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(G211gat), .B(G218gat), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G204gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G197gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT96), .ZN(new_n340_));
  INV_X1    g139(.A(new_n338_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(KEYINPUT96), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n334_), .B(new_n336_), .C1(new_n344_), .C2(KEYINPUT21), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n342_), .B1(new_n339_), .B2(KEYINPUT96), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT97), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT21), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n335_), .B1(new_n346_), .B2(KEYINPUT97), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n345_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n330_), .B1(new_n331_), .B2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n313_), .A2(new_n314_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT93), .B1(new_n319_), .B2(new_n323_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT29), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n330_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n351_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n329_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G22gat), .B(G50gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n355_), .B1(new_n325_), .B2(KEYINPUT29), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n328_), .B(new_n326_), .C1(new_n362_), .C2(new_n351_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n358_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n361_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n265_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT103), .ZN(new_n368_));
  INV_X1    g167(.A(new_n260_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n315_), .B2(new_n324_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT101), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT100), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n313_), .A2(new_n260_), .ZN(new_n374_));
  NOR4_X1   g173(.A1(new_n370_), .A2(new_n371_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n325_), .B2(new_n260_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n373_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT101), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n260_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n374_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n379_), .A2(KEYINPUT99), .A3(KEYINPUT4), .A4(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n370_), .A2(new_n382_), .A3(new_n374_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n382_), .B(new_n260_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT99), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n381_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n387_));
  AOI211_X1 g186(.A(new_n375_), .B(new_n378_), .C1(new_n387_), .C2(new_n373_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  INV_X1    g188(.A(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n368_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n388_), .A2(new_n394_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n387_), .A2(new_n373_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n375_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n378_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(KEYINPUT103), .A3(new_n393_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(new_n396_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT19), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n242_), .B2(new_n350_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n204_), .A2(new_n206_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n209_), .A2(new_n211_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n227_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT98), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n218_), .B(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n238_), .B(new_n410_), .C1(new_n219_), .C2(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT22), .B(G169gat), .Z(new_n414_));
  INV_X1    g213(.A(new_n225_), .ZN(new_n415_));
  OAI221_X1 g214(.A(new_n217_), .B1(new_n414_), .B2(G176gat), .C1(new_n415_), .C2(new_n240_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n350_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n405_), .B1(new_n407_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT97), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n344_), .A2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n421_), .A2(KEYINPUT21), .A3(new_n335_), .A4(new_n347_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n229_), .A2(new_n422_), .A3(new_n345_), .A4(new_n241_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n350_), .A2(new_n417_), .ZN(new_n424_));
  AND4_X1   g223(.A1(KEYINPUT20), .A2(new_n423_), .A3(new_n424_), .A4(new_n405_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n419_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n404_), .B1(new_n407_), .B2(new_n418_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n423_), .A2(new_n424_), .A3(KEYINPUT20), .A4(new_n404_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n426_), .B1(new_n430_), .B2(KEYINPUT102), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(G92gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT18), .B(G64gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n433_), .B(new_n434_), .Z(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT32), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n430_), .A2(new_n437_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n431_), .A2(new_n437_), .B1(new_n438_), .B2(KEYINPUT102), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n402_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n396_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n388_), .A2(KEYINPUT33), .A3(new_n394_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n435_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n407_), .A2(new_n418_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n428_), .B(new_n444_), .C1(new_n445_), .C2(new_n404_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n435_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n387_), .A2(new_n377_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n376_), .A2(new_n373_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n393_), .A3(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n442_), .A2(new_n443_), .A3(new_n448_), .A4(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n367_), .B1(new_n440_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n265_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n444_), .B1(new_n419_), .B2(new_n425_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n447_), .A2(new_n455_), .A3(KEYINPUT27), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT27), .B1(new_n446_), .B2(new_n447_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT104), .B1(new_n366_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n358_), .A2(new_n363_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n361_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n358_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n463_));
  AND4_X1   g262(.A1(KEYINPUT104), .A2(new_n462_), .A3(new_n458_), .A4(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n454_), .B1(new_n459_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n366_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(new_n265_), .A3(new_n458_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n402_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n453_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G43gat), .B(G50gat), .Z(new_n470_));
  XNOR2_X1  g269(.A(G29gat), .B(G36gat), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n471_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n474_), .B(KEYINPUT15), .Z(new_n475_));
  XNOR2_X1  g274(.A(G85gat), .B(G92gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT9), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT10), .B(G99gat), .Z(new_n479_));
  INV_X1    g278(.A(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482_));
  INV_X1    g281(.A(G99gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n480_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n477_), .A2(G85gat), .A3(G92gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n478_), .A2(new_n481_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n476_), .A2(KEYINPUT65), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n483_), .A2(new_n480_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT64), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n490_), .B(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n484_), .B(new_n485_), .C1(KEYINPUT64), .C2(new_n491_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n489_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n495_), .A2(KEYINPUT8), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n497_), .B(new_n489_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n488_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G232gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT34), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT35), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n475_), .A2(new_n500_), .B1(KEYINPUT70), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n488_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n495_), .A2(KEYINPUT8), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(new_n498_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n505_), .B(new_n509_), .C1(KEYINPUT35), .C2(new_n502_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n504_), .A2(KEYINPUT70), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G190gat), .B(G218gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G162gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT69), .B(G134gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT36), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(KEYINPUT71), .A2(KEYINPUT72), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(KEYINPUT37), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT71), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(new_n518_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n512_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n516_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n518_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(KEYINPUT72), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530_));
  INV_X1    g329(.A(G1gat), .ZN(new_n531_));
  INV_X1    g330(.A(G8gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT14), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G1gat), .B(G8gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT73), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n536_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n542_));
  XOR2_X1   g341(.A(G71gat), .B(G78gat), .Z(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n542_), .A2(new_n543_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n539_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT76), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G127gat), .B(G155gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G211gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT16), .B(G183gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT17), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT74), .B(KEYINPUT17), .Z(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT75), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(new_n547_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n526_), .A2(new_n529_), .A3(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT77), .Z(new_n562_));
  AND2_X1   g361(.A1(new_n469_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT68), .ZN(new_n565_));
  INV_X1    g364(.A(new_n546_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT12), .B1(new_n500_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n508_), .A2(new_n568_), .A3(new_n546_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n488_), .B(new_n546_), .C1(new_n496_), .C2(new_n499_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT66), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT66), .ZN(new_n574_));
  INV_X1    g373(.A(new_n572_), .ZN(new_n575_));
  AOI211_X1 g374(.A(new_n574_), .B(new_n575_), .C1(new_n508_), .C2(new_n546_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n570_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n571_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n508_), .A2(new_n546_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n575_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(G204gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT5), .B(G176gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  OR2_X1    g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT67), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(new_n585_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n581_), .A2(KEYINPUT67), .A3(new_n585_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n565_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n564_), .A2(KEYINPUT68), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n592_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n536_), .B(new_n474_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n536_), .A2(new_n474_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n475_), .B2(new_n536_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600_));
  MUX2_X1   g399(.A(new_n597_), .B(new_n599_), .S(new_n600_), .Z(new_n601_));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n601_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n596_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n563_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(new_n531_), .A3(new_n402_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT38), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n469_), .A2(new_n528_), .A3(new_n607_), .A4(new_n560_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n402_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(G1324gat));
  AND2_X1   g414(.A1(new_n469_), .A2(new_n528_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n458_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n616_), .A2(new_n617_), .A3(new_n607_), .A4(new_n560_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT105), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(G8gat), .A3(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n609_), .A2(new_n532_), .A3(new_n617_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n622_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n618_), .A2(G8gat), .A3(new_n620_), .A4(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n623_), .A2(KEYINPUT40), .A3(new_n624_), .A4(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1325gat));
  OAI21_X1  g430(.A(G15gat), .B1(new_n612_), .B2(new_n265_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n265_), .A2(G15gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n608_), .B2(new_n635_), .ZN(G1326gat));
  OR3_X1    g435(.A1(new_n608_), .A2(G22gat), .A3(new_n366_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G22gat), .B1(new_n612_), .B2(new_n366_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT107), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(KEYINPUT107), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n640_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n637_), .B1(new_n642_), .B2(new_n643_), .ZN(G1327gat));
  INV_X1    g443(.A(G29gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n526_), .A2(new_n529_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n646_), .B1(new_n453_), .B2(new_n468_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT43), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n649_), .B(new_n646_), .C1(new_n453_), .C2(new_n468_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n596_), .A2(new_n606_), .A3(new_n560_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n651_), .A2(KEYINPUT108), .A3(new_n652_), .A4(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n657_));
  OAI21_X1  g456(.A(new_n654_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n645_), .B1(new_n658_), .B2(new_n402_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n528_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n653_), .B(new_n660_), .C1(new_n468_), .C2(new_n453_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n661_), .A2(G29gat), .A3(new_n613_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT109), .B1(new_n659_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT109), .ZN(new_n664_));
  INV_X1    g463(.A(new_n662_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n657_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n613_), .B1(new_n667_), .B2(new_n654_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n664_), .B(new_n665_), .C1(new_n668_), .C2(new_n645_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n663_), .A2(new_n669_), .ZN(G1328gat));
  XNOR2_X1  g469(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n652_), .A2(KEYINPUT108), .ZN(new_n672_));
  AOI211_X1 g471(.A(new_n655_), .B(new_n672_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n617_), .B1(new_n666_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G36gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n661_), .ZN(new_n676_));
  INV_X1    g475(.A(G36gat), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(KEYINPUT45), .A3(new_n677_), .A4(new_n617_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n469_), .A2(new_n677_), .A3(new_n660_), .A4(new_n653_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(new_n458_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n671_), .B1(new_n675_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n671_), .ZN(new_n685_));
  AOI211_X1 g484(.A(new_n685_), .B(new_n682_), .C1(new_n674_), .C2(G36gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1329gat));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n454_), .B1(new_n666_), .B2(new_n673_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G43gat), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n661_), .A2(G43gat), .A3(new_n265_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n688_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT47), .B(new_n691_), .C1(new_n689_), .C2(G43gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1330gat));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n658_), .A2(new_n696_), .A3(new_n466_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n466_), .B1(new_n666_), .B2(new_n673_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT111), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n699_), .A3(G50gat), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n366_), .A2(G50gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n661_), .B2(new_n701_), .ZN(G1331gat));
  NOR2_X1   g501(.A1(new_n595_), .A2(new_n605_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n616_), .A2(new_n560_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n613_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n563_), .A2(new_n703_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT112), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n563_), .A2(KEYINPUT112), .A3(new_n703_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n402_), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n705_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT113), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(KEYINPUT113), .A3(new_n705_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n706_), .B1(new_n714_), .B2(new_n715_), .ZN(G1332gat));
  AND2_X1   g515(.A1(new_n709_), .A2(new_n710_), .ZN(new_n717_));
  INV_X1    g516(.A(G64gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n617_), .ZN(new_n719_));
  AND4_X1   g518(.A1(new_n617_), .A2(new_n616_), .A3(new_n560_), .A4(new_n703_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT114), .B1(new_n720_), .B2(new_n718_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n723_), .B(G64gat), .C1(new_n704_), .C2(new_n458_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n721_), .A2(new_n722_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n722_), .B1(new_n721_), .B2(new_n724_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n719_), .B1(new_n725_), .B2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n704_), .B2(new_n265_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n717_), .A2(new_n731_), .A3(new_n454_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n704_), .B2(new_n366_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  INV_X1    g534(.A(G78gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n717_), .A2(new_n736_), .A3(new_n466_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1335gat));
  AND2_X1   g537(.A1(new_n469_), .A2(new_n660_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n703_), .A2(new_n559_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n402_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n740_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n613_), .A2(new_n390_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(G1336gat));
  AOI21_X1  g546(.A(G92gat), .B1(new_n743_), .B2(new_n617_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n617_), .A2(G92gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n745_), .B2(new_n749_), .ZN(G1337gat));
  NAND3_X1  g549(.A1(new_n743_), .A2(new_n479_), .A3(new_n454_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n745_), .A2(new_n454_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n483_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT51), .ZN(G1338gat));
  AND4_X1   g553(.A1(new_n480_), .A2(new_n739_), .A3(new_n466_), .A4(new_n741_), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n366_), .B(new_n740_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT52), .B1(new_n756_), .B2(new_n480_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n745_), .A2(new_n466_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n755_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n762_), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n764_), .B(new_n755_), .C1(new_n757_), .C2(new_n760_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1339gat));
  OR2_X1    g565(.A1(new_n459_), .A2(new_n464_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n402_), .A3(new_n454_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n576_), .A2(new_n573_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n569_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n568_), .B1(new_n508_), .B2(new_n546_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n575_), .B1(new_n773_), .B2(new_n578_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n570_), .B(KEYINPUT55), .C1(new_n573_), .C2(new_n576_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n585_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  MUX2_X1   g581(.A(new_n599_), .B(new_n597_), .S(new_n600_), .Z(new_n783_));
  MUX2_X1   g582(.A(new_n601_), .B(new_n783_), .S(new_n604_), .Z(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n586_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n782_), .A2(KEYINPUT58), .A3(new_n586_), .A4(new_n784_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n646_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n780_), .A2(new_n791_), .A3(new_n781_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n777_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n585_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n605_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n794_), .A3(new_n586_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n589_), .A2(new_n590_), .A3(new_n784_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n790_), .B1(new_n797_), .B2(new_n528_), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT57), .B(new_n660_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n789_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT118), .B(new_n789_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n559_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n561_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n595_), .A2(new_n805_), .A3(new_n806_), .A4(new_n606_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n593_), .A2(new_n606_), .A3(new_n594_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT54), .B1(new_n808_), .B2(new_n561_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n768_), .B1(new_n804_), .B2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(G113gat), .B1(new_n811_), .B2(new_n605_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n813_), .B(new_n768_), .C1(new_n804_), .C2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n800_), .A2(new_n559_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n815_), .A2(new_n810_), .B1(new_n816_), .B2(new_n768_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n768_), .A2(new_n816_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT59), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n814_), .A2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(new_n605_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n812_), .B1(new_n821_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n595_), .B2(G120gat), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n811_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n823_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n596_), .B1(new_n814_), .B2(new_n819_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT120), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n829_), .B(new_n596_), .C1(new_n814_), .C2(new_n819_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n825_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n826_), .B1(new_n831_), .B2(new_n832_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n811_), .B2(new_n560_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n820_), .A2(new_n560_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g635(.A(G134gat), .B1(new_n811_), .B2(new_n660_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n820_), .A2(new_n646_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g638(.A1(new_n613_), .A2(new_n467_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT121), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n804_), .B2(new_n810_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n605_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n596_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n560_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n847_), .A2(G155gat), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(G155gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n850_), .B(new_n852_), .ZN(G1346gat));
  AOI21_X1  g652(.A(G162gat), .B1(new_n842_), .B2(new_n660_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n646_), .A2(G162gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n842_), .B2(new_n855_), .ZN(G1347gat));
  NAND2_X1  g655(.A1(new_n613_), .A2(new_n617_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n366_), .A3(new_n454_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n810_), .B2(new_n815_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n605_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G169gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT123), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n864_), .A3(G169gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n863_), .A2(KEYINPUT62), .A3(new_n865_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n868_), .B(new_n869_), .C1(new_n414_), .C2(new_n861_), .ZN(G1348gat));
  AOI21_X1  g669(.A(G176gat), .B1(new_n860_), .B2(new_n596_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n859_), .B1(new_n804_), .B2(new_n810_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n596_), .A2(G176gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1349gat));
  INV_X1    g673(.A(new_n860_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n875_), .A2(new_n409_), .A3(new_n559_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G183gat), .B1(new_n872_), .B2(new_n560_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1350gat));
  INV_X1    g677(.A(new_n646_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G190gat), .B1(new_n875_), .B2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n860_), .A2(new_n660_), .A3(new_n408_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1351gat));
  AOI211_X1 g681(.A(new_n366_), .B(new_n454_), .C1(new_n804_), .C2(new_n810_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n858_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G197gat), .B1(new_n885_), .B2(new_n605_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n883_), .A2(G197gat), .A3(new_n605_), .A4(new_n858_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(KEYINPUT124), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(KEYINPUT124), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n886_), .A2(new_n888_), .A3(new_n889_), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n885_), .A2(new_n596_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT125), .B(G204gat), .Z(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(new_n893_), .ZN(G1353gat));
  NOR2_X1   g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  AND2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n884_), .A2(new_n559_), .A3(new_n895_), .A4(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n884_), .B2(new_n559_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT126), .B(new_n895_), .C1(new_n884_), .C2(new_n559_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  OAI21_X1  g701(.A(G218gat), .B1(new_n884_), .B2(new_n879_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n528_), .A2(G218gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n883_), .A2(new_n858_), .A3(new_n905_), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n903_), .A2(new_n904_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n904_), .B1(new_n903_), .B2(new_n906_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1355gat));
endmodule


