//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n978_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n985_, new_n986_, new_n987_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n216_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT10), .B(G99gat), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT65), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT10), .B(G99gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n222_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n229_));
  INV_X1    g028(.A(G85gat), .ZN(new_n230_));
  INV_X1    g029(.A(G92gat), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT9), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n212_), .A2(new_n213_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OAI22_X1  g033(.A1(new_n219_), .A2(new_n220_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G29gat), .B(G36gat), .Z(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(KEYINPUT73), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G29gat), .B(G36gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT73), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(G43gat), .B1(new_n237_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(KEYINPUT73), .ZN(new_n242_));
  INV_X1    g041(.A(G43gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n239_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n241_), .A2(G50gat), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(G50gat), .B1(new_n241_), .B2(new_n245_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT15), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G50gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n245_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n243_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n241_), .A2(G50gat), .A3(new_n245_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT15), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n235_), .B1(new_n249_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n254_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(new_n235_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT34), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT35), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n228_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n234_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n220_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n265_), .A2(new_n266_), .B1(new_n267_), .B2(new_n218_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n248_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n253_), .A2(KEYINPUT15), .A3(new_n254_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n264_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n262_), .A2(KEYINPUT35), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n260_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n269_), .A2(new_n270_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n258_), .B1(new_n277_), .B2(new_n235_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n256_), .A2(KEYINPUT74), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(new_n264_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n205_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n273_), .A2(new_n260_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n204_), .B(KEYINPUT36), .Z(new_n283_));
  AOI21_X1  g082(.A(new_n274_), .B1(new_n279_), .B2(new_n264_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n282_), .B(new_n283_), .C1(new_n284_), .C2(new_n260_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT37), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n281_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n263_), .B1(new_n256_), .B2(KEYINPUT74), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n278_), .B1(new_n288_), .B2(new_n274_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n283_), .B(KEYINPUT75), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n282_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n281_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT76), .B1(new_n287_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n290_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n276_), .A2(new_n280_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n205_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n289_), .B2(new_n282_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT37), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n281_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n293_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G127gat), .B(G155gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT16), .ZN(new_n304_));
  INV_X1    g103(.A(G183gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(G211gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT17), .ZN(new_n308_));
  INV_X1    g107(.A(G1gat), .ZN(new_n309_));
  INV_X1    g108(.A(G8gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT14), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT77), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n313_), .B(KEYINPUT14), .C1(new_n309_), .C2(new_n310_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G15gat), .B(G22gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G1gat), .B(G8gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G231gat), .A2(G233gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(KEYINPUT78), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n318_), .B(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G57gat), .B(G64gat), .Z(new_n322_));
  INV_X1    g121(.A(KEYINPUT11), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G71gat), .B(G78gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(G57gat), .B(G64gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(KEYINPUT11), .B2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n328_), .A2(KEYINPUT67), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n322_), .A2(new_n323_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n330_), .B1(new_n331_), .B2(new_n326_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n325_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(KEYINPUT67), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n330_), .A3(new_n326_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n324_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n321_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n321_), .A2(new_n337_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n308_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT80), .Z(new_n341_));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n333_), .A2(KEYINPUT69), .A3(new_n336_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(new_n321_), .Z(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n346_), .A2(new_n307_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n341_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n302_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(KEYINPUT81), .Z(new_n351_));
  NAND2_X1  g150(.A1(G230gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT64), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n337_), .A2(new_n268_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT68), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n235_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n343_), .A2(new_n344_), .A3(KEYINPUT12), .A4(new_n235_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n337_), .B2(new_n268_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT70), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT12), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n356_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n359_), .B(new_n360_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n366_));
  XNOR2_X1  g165(.A(G120gat), .B(G148gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G176gat), .B(G204gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  NAND3_X1  g169(.A1(new_n358_), .A2(new_n365_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n358_), .B2(new_n365_), .ZN(new_n373_));
  AND2_X1   g172(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n374_));
  OR3_X1    g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n376_));
  OAI22_X1  g175(.A1(new_n372_), .A2(new_n373_), .B1(new_n376_), .B2(new_n374_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n351_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT18), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G64gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G92gat), .ZN(new_n384_));
  INV_X1    g183(.A(G64gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n382_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n231_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT19), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT23), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT23), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(G183gat), .A3(G190gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n393_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n305_), .A2(KEYINPUT82), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G183gat), .ZN(new_n400_));
  INV_X1    g199(.A(G190gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n394_), .A2(KEYINPUT86), .A3(G183gat), .A4(G190gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n397_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G169gat), .ZN(new_n405_));
  INV_X1    g204(.A(G176gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n409_));
  NAND2_X1  g208(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n410_));
  AOI21_X1  g209(.A(G176gat), .B1(new_n410_), .B2(G169gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n405_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(G169gat), .ZN(new_n414_));
  AND4_X1   g213(.A1(new_n409_), .A2(new_n414_), .A3(new_n412_), .A4(new_n406_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n404_), .B(new_n408_), .C1(new_n413_), .C2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT83), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n393_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n392_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n395_), .A3(new_n419_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT24), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(G169gat), .B2(G176gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G169gat), .A2(G176gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n421_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n398_), .A2(new_n400_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(KEYINPUT25), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT26), .B(G190gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n420_), .B(new_n426_), .C1(new_n429_), .C2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n416_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G197gat), .B(G204gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(G211gat), .B(G218gat), .Z(new_n435_));
  INV_X1    g234(.A(KEYINPUT21), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G211gat), .B(G218gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT21), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n434_), .A3(KEYINPUT21), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT90), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT90), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n433_), .A2(new_n445_), .A3(new_n442_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n444_), .A2(KEYINPUT20), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n421_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n397_), .A2(new_n403_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n423_), .A2(new_n425_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n397_), .A2(KEYINPUT89), .A3(new_n403_), .A4(new_n448_), .ZN(new_n453_));
  OR2_X1    g252(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT88), .ZN(new_n455_));
  NAND2_X1  g254(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT88), .B1(new_n458_), .B2(new_n427_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n430_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .A4(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n420_), .B1(G183gat), .B2(G190gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT22), .B(G169gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n407_), .B1(new_n464_), .B2(new_n406_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT94), .ZN(new_n468_));
  INV_X1    g267(.A(new_n442_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n470_), .A3(new_n466_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n391_), .B1(new_n447_), .B2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n469_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT20), .B1(new_n433_), .B2(new_n442_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n390_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n388_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n462_), .A2(new_n466_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n390_), .B1(new_n478_), .B2(new_n469_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n443_), .B2(KEYINPUT90), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n446_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n388_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n390_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n477_), .A2(KEYINPUT27), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G155gat), .B(G162gat), .ZN(new_n487_));
  INV_X1    g286(.A(G141gat), .ZN(new_n488_));
  INV_X1    g287(.A(G148gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT3), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT3), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(G141gat), .B2(G148gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n487_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(G155gat), .A2(G162gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G155gat), .A2(G162gat), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT1), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n488_), .A2(new_n489_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G141gat), .A2(G148gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT29), .B1(new_n497_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n442_), .A2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(G228gat), .A2(G233gat), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n508_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n497_), .A2(new_n505_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G22gat), .B(G50gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT28), .ZN(new_n517_));
  XOR2_X1   g316(.A(G78gat), .B(G106gat), .Z(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OR3_X1    g319(.A1(new_n514_), .A2(new_n515_), .A3(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT27), .ZN(new_n524_));
  INV_X1    g323(.A(new_n485_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n483_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n486_), .A2(new_n523_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G1gat), .B(G29gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT0), .ZN(new_n531_));
  INV_X1    g330(.A(G57gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G85gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G134gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(G127gat), .ZN(new_n537_));
  INV_X1    g336(.A(G127gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(G134gat), .ZN(new_n539_));
  INV_X1    g338(.A(G120gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(G113gat), .ZN(new_n541_));
  INV_X1    g340(.A(G113gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G120gat), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n537_), .A2(new_n539_), .A3(new_n541_), .A4(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n537_), .A2(new_n539_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n544_), .B(new_n547_), .C1(new_n497_), .C2(new_n505_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n487_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n490_), .A2(new_n492_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n495_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n549_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n501_), .A2(new_n502_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n555_), .B(new_n503_), .C1(KEYINPUT1), .C2(new_n487_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(new_n544_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n548_), .A2(new_n558_), .A3(KEYINPUT91), .ZN(new_n559_));
  INV_X1    g358(.A(new_n557_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n560_), .B(new_n561_), .C1(new_n497_), .C2(new_n505_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(KEYINPUT4), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT4), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n548_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G225gat), .A2(G233gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n559_), .A2(new_n562_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT92), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n568_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n535_), .B1(new_n570_), .B2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n569_), .A2(new_n573_), .A3(new_n534_), .A4(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G15gat), .B(G43gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT31), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n433_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n416_), .A2(KEYINPUT30), .A3(new_n432_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G227gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT87), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G71gat), .B(G99gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n587_), .A2(new_n592_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n557_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n557_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n583_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n598_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n582_), .A3(new_n596_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n580_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n529_), .A2(KEYINPUT97), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n601_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n580_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n604_), .B1(new_n607_), .B2(new_n528_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n521_), .A2(new_n522_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n472_), .A2(new_n446_), .A3(new_n481_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n476_), .B1(new_n613_), .B2(new_n390_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n384_), .A2(new_n387_), .A3(KEYINPUT32), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  OAI211_X1 g416(.A(KEYINPUT95), .B(new_n617_), .C1(new_n473_), .C2(new_n476_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n444_), .A2(KEYINPUT20), .A3(new_n446_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n391_), .B1(new_n467_), .B2(new_n442_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n484_), .B(new_n615_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT93), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n482_), .A2(KEYINPUT93), .A3(new_n615_), .A4(new_n484_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n578_), .A2(new_n579_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n619_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n579_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n574_), .B(KEYINPUT92), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n630_), .A2(KEYINPUT33), .A3(new_n534_), .A4(new_n569_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n566_), .A2(new_n567_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n571_), .A2(new_n568_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n535_), .A3(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n629_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n525_), .A2(new_n526_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n611_), .B1(new_n627_), .B2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n606_), .A2(new_n486_), .A3(new_n611_), .A4(new_n527_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n610_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT96), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n643_), .B(new_n610_), .C1(new_n638_), .C2(new_n640_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n609_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n318_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n257_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n277_), .A2(new_n646_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n257_), .B(new_n646_), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n650_), .A2(new_n651_), .B1(new_n652_), .B2(new_n649_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G113gat), .B(G141gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(new_n405_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(G197gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n653_), .B(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT98), .B1(new_n645_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n603_), .A2(new_n608_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n644_), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n619_), .A2(new_n626_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n639_), .B1(new_n662_), .B2(new_n611_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n643_), .B1(new_n663_), .B2(new_n610_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n661_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n657_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n659_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n380_), .A2(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n669_), .A2(G1gat), .A3(new_n606_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n349_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n281_), .A2(new_n285_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n645_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n379_), .A2(new_n658_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT100), .ZN(new_n679_));
  OAI21_X1  g478(.A(G1gat), .B1(new_n679_), .B2(new_n606_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n672_), .A2(new_n680_), .ZN(G1324gat));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n477_), .A2(KEYINPUT27), .A3(new_n485_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n526_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT27), .B1(new_n684_), .B2(new_n485_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n676_), .A2(new_n677_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT39), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(new_n689_), .A3(G8gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(G8gat), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n380_), .A2(new_n310_), .A3(new_n687_), .A4(new_n668_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n682_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n697_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(KEYINPUT40), .A3(new_n695_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1325gat));
  OR3_X1    g500(.A1(new_n669_), .A2(G15gat), .A3(new_n610_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G15gat), .B1(new_n679_), .B2(new_n610_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n703_), .A2(new_n704_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1326gat));
  OAI21_X1  g506(.A(G22gat), .B1(new_n679_), .B2(new_n523_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT42), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n523_), .A2(G22gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n669_), .B2(new_n710_), .ZN(G1327gat));
  NOR2_X1   g510(.A1(new_n673_), .A2(new_n674_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n378_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n659_), .B2(new_n667_), .ZN(new_n714_));
  INV_X1    g513(.A(G29gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n580_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n677_), .A2(new_n349_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n293_), .A2(new_n301_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n645_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n665_), .A2(new_n720_), .A3(new_n302_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n717_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT44), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n580_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n717_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n645_), .A2(KEYINPUT43), .A3(new_n718_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n720_), .B1(new_n665_), .B2(new_n302_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n728_), .B2(KEYINPUT102), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT102), .B(new_n717_), .C1(new_n719_), .C2(new_n721_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n729_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n722_), .B2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT103), .B1(new_n736_), .B2(new_n730_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n724_), .B1(new_n733_), .B2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738_), .B2(KEYINPUT104), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n740_));
  AOI211_X1 g539(.A(new_n740_), .B(new_n724_), .C1(new_n733_), .C2(new_n737_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n716_), .B1(new_n739_), .B2(new_n741_), .ZN(G1328gat));
  NOR2_X1   g541(.A1(new_n686_), .A2(G36gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n714_), .A2(new_n743_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(KEYINPUT45), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(KEYINPUT45), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n723_), .A2(new_n687_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n733_), .B2(new_n737_), .ZN(new_n750_));
  INV_X1    g549(.A(G36gat), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n748_), .B(KEYINPUT46), .C1(new_n750_), .C2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n749_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n732_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n736_), .A2(KEYINPUT103), .A3(new_n730_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n747_), .B1(new_n756_), .B2(G36gat), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n752_), .B1(new_n757_), .B2(new_n758_), .ZN(G1329gat));
  NAND3_X1  g558(.A1(new_n723_), .A2(G43gat), .A3(new_n605_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n733_), .B2(new_n737_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G43gat), .B1(new_n714_), .B2(new_n605_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(KEYINPUT106), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(KEYINPUT106), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OR3_X1    g564(.A1(new_n761_), .A2(new_n765_), .A3(KEYINPUT47), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT47), .B1(new_n761_), .B2(new_n765_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1330gat));
  AOI21_X1  g567(.A(G50gat), .B1(new_n714_), .B2(new_n611_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n733_), .A2(new_n737_), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n250_), .B(new_n523_), .C1(new_n722_), .C2(KEYINPUT44), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n770_), .B2(new_n771_), .ZN(G1331gat));
  NOR2_X1   g571(.A1(new_n378_), .A2(new_n657_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n676_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G57gat), .B1(new_n774_), .B2(new_n606_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n773_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n351_), .A2(new_n645_), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n580_), .A2(new_n532_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT107), .Z(G1332gat));
  OAI21_X1  g580(.A(G64gat), .B1(new_n774_), .B2(new_n686_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT48), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n777_), .A2(new_n385_), .A3(new_n687_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1333gat));
  OAI21_X1  g584(.A(G71gat), .B1(new_n774_), .B2(new_n610_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT49), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n610_), .A2(G71gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n778_), .B2(new_n788_), .ZN(G1334gat));
  OAI21_X1  g588(.A(G78gat), .B1(new_n774_), .B2(new_n523_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT50), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n523_), .A2(G78gat), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT108), .Z(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n778_), .B2(new_n793_), .ZN(G1335gat));
  NOR2_X1   g593(.A1(new_n726_), .A2(new_n727_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n795_), .A2(KEYINPUT110), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(KEYINPUT110), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n776_), .A2(new_n673_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799_), .B2(new_n606_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n665_), .A2(new_n712_), .A3(new_n773_), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT109), .Z(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(new_n230_), .A3(new_n580_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n803_), .ZN(G1336gat));
  OAI21_X1  g603(.A(G92gat), .B1(new_n799_), .B2(new_n686_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(new_n231_), .A3(new_n687_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT111), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n809_), .A3(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1337gat));
  NAND4_X1  g610(.A1(new_n796_), .A2(new_n797_), .A3(new_n605_), .A4(new_n798_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G99gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n610_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT112), .B1(new_n802_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1338gat));
  NAND2_X1  g617(.A1(new_n798_), .A2(new_n611_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G106gat), .B1(new_n795_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT52), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n802_), .A2(new_n221_), .A3(new_n611_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n365_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n356_), .A2(new_n362_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT70), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n356_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n831_), .A2(KEYINPUT55), .A3(new_n359_), .A4(new_n360_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n827_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n359_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n353_), .B1(new_n834_), .B2(new_n355_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT68), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n354_), .B(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n831_), .A3(new_n359_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(KEYINPUT114), .A3(new_n353_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n833_), .B1(new_n837_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n825_), .B1(new_n842_), .B2(new_n370_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n827_), .A2(new_n832_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n835_), .A2(new_n836_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT114), .B1(new_n840_), .B2(new_n353_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n370_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(KEYINPUT56), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n843_), .A2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n651_), .B(new_n649_), .C1(new_n646_), .C2(new_n257_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n656_), .B1(new_n652_), .B2(new_n648_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n653_), .A2(new_n656_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n371_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT116), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n850_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n718_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n850_), .A2(KEYINPUT58), .A3(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n657_), .A2(new_n371_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n843_), .B2(new_n849_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n853_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT115), .B(new_n853_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(KEYINPUT57), .B(new_n674_), .C1(new_n862_), .C2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n674_), .B1(new_n862_), .B2(new_n867_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n860_), .A2(new_n868_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n673_), .B1(new_n872_), .B2(KEYINPUT117), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n858_), .A2(new_n859_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n868_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n350_), .A2(new_n658_), .A3(new_n378_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT54), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n877_), .A2(KEYINPUT54), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n873_), .A2(new_n876_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n610_), .A2(new_n606_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n529_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n542_), .A3(new_n657_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n872_), .A2(KEYINPUT117), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n349_), .A3(new_n876_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n877_), .B(KEYINPUT54), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n882_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n886_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n886_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n868_), .B1(new_n874_), .B2(KEYINPUT118), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n860_), .A2(KEYINPUT118), .A3(new_n871_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n349_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n896_), .B2(new_n889_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n885_), .B1(new_n892_), .B2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT59), .B1(new_n880_), .B2(new_n882_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n897_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n900_), .A3(KEYINPUT119), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n658_), .B1(new_n898_), .B2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n884_), .B1(new_n902_), .B2(new_n542_), .ZN(G1340gat));
  OAI21_X1  g702(.A(new_n540_), .B1(new_n378_), .B2(KEYINPUT60), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n883_), .B(new_n904_), .C1(KEYINPUT60), .C2(new_n540_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n892_), .A2(new_n378_), .A3(new_n897_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n540_), .ZN(G1341gat));
  NAND3_X1  g706(.A1(new_n883_), .A2(new_n538_), .A3(new_n673_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n349_), .B1(new_n898_), .B2(new_n901_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n538_), .ZN(G1342gat));
  INV_X1    g709(.A(new_n674_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n883_), .A2(new_n536_), .A3(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n718_), .B1(new_n898_), .B2(new_n901_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n536_), .ZN(G1343gat));
  NOR4_X1   g713(.A1(new_n687_), .A2(new_n606_), .A3(new_n523_), .A4(new_n605_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n890_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT120), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n890_), .A2(new_n918_), .A3(new_n915_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n658_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT121), .B(G141gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1344gat));
  AOI21_X1  g721(.A(new_n378_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n489_), .ZN(G1345gat));
  AOI21_X1  g723(.A(new_n349_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT61), .B(G155gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT122), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n925_), .B(new_n927_), .ZN(G1346gat));
  NAND2_X1  g727(.A1(new_n917_), .A2(new_n919_), .ZN(new_n929_));
  INV_X1    g728(.A(G162gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(new_n930_), .A3(new_n911_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n718_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n930_), .ZN(G1347gat));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n686_), .A2(new_n607_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n611_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n896_), .B2(new_n889_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n939_), .A2(new_n657_), .A3(new_n464_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n405_), .B1(new_n939_), .B2(new_n657_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(KEYINPUT62), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n943_));
  AOI211_X1 g742(.A(new_n943_), .B(new_n405_), .C1(new_n939_), .C2(new_n657_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n934_), .B1(new_n942_), .B2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n896_), .A2(new_n889_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n946_), .A2(new_n657_), .A3(new_n937_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(G169gat), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n943_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n941_), .A2(KEYINPUT62), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n949_), .A2(new_n950_), .A3(KEYINPUT123), .A4(new_n940_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n945_), .A2(new_n951_), .ZN(G1348gat));
  AOI21_X1  g751(.A(G176gat), .B1(new_n939_), .B2(new_n379_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n379_), .A2(G176gat), .A3(new_n935_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n880_), .A2(new_n611_), .A3(new_n954_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n953_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n956_), .B(new_n957_), .ZN(G1349gat));
  NOR2_X1   g757(.A1(new_n880_), .A2(new_n611_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n936_), .A2(new_n349_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(KEYINPUT125), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n959_), .A2(new_n963_), .A3(new_n960_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n428_), .B1(new_n962_), .B2(new_n964_), .ZN(new_n965_));
  INV_X1    g764(.A(new_n939_), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n966_), .A2(new_n460_), .A3(new_n349_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n965_), .A2(new_n967_), .ZN(G1350gat));
  OAI21_X1  g767(.A(G190gat), .B1(new_n966_), .B2(new_n718_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n939_), .A2(new_n430_), .A3(new_n911_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1351gat));
  NOR3_X1   g770(.A1(new_n605_), .A2(new_n523_), .A3(new_n580_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n972_), .A2(KEYINPUT126), .ZN(new_n973_));
  AND2_X1   g772(.A1(new_n972_), .A2(KEYINPUT126), .ZN(new_n974_));
  NOR4_X1   g773(.A1(new_n880_), .A2(new_n686_), .A3(new_n973_), .A4(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(new_n657_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n379_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g778(.A1(new_n975_), .A2(new_n673_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(KEYINPUT63), .B(G211gat), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n980_), .A2(new_n981_), .ZN(new_n982_));
  NOR2_X1   g781(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n982_), .B1(new_n980_), .B2(new_n983_), .ZN(G1354gat));
  NAND2_X1  g783(.A1(new_n975_), .A2(new_n911_), .ZN(new_n985_));
  XOR2_X1   g784(.A(KEYINPUT127), .B(G218gat), .Z(new_n986_));
  NOR2_X1   g785(.A1(new_n718_), .A2(new_n986_), .ZN(new_n987_));
  AOI22_X1  g786(.A1(new_n985_), .A2(new_n986_), .B1(new_n975_), .B2(new_n987_), .ZN(G1355gat));
endmodule


