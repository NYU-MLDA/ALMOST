//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  OR2_X1    g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT24), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n219_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT77), .B(G190gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n227_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n226_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G183gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n234_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n235_), .A2(new_n219_), .B1(G169gat), .B2(G176gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n220_), .A2(KEYINPUT22), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n237_), .A2(KEYINPUT78), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(KEYINPUT78), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT22), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G169gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n238_), .A2(new_n239_), .A3(new_n221_), .A4(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n214_), .A2(new_n233_), .A3(new_n243_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n217_), .B(new_n218_), .C1(G183gat), .C2(G190gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n241_), .A3(new_n221_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n224_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT26), .B(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n227_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n226_), .A2(KEYINPUT91), .A3(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n250_), .A2(new_n219_), .A3(new_n223_), .A4(new_n225_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT91), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n248_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(KEYINPUT20), .B(new_n244_), .C1(new_n255_), .C2(new_n214_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G226gat), .A2(G233gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT19), .Z(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G8gat), .B(G36gat), .Z(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT18), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G64gat), .B(G92gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n255_), .A2(new_n214_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(KEYINPUT20), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n233_), .A2(new_n243_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(new_n213_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n260_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n264_), .B1(new_n260_), .B2(new_n269_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n203_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n256_), .A2(new_n259_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n203_), .B1(new_n273_), .B2(new_n264_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n264_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n256_), .A2(new_n259_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT20), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n267_), .B2(new_n213_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n214_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n258_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n275_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n274_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(G15gat), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G71gat), .B(G99gat), .Z(new_n286_));
  INV_X1    g085(.A(G43gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G71gat), .B(G99gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G43gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT30), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n293_), .A3(new_n290_), .ZN(new_n294_));
  AND4_X1   g093(.A1(new_n233_), .A2(new_n243_), .A3(new_n292_), .A4(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n233_), .A2(new_n243_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n285_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT80), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n292_), .A2(new_n294_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n267_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n233_), .A2(new_n243_), .A3(new_n292_), .A4(new_n294_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n284_), .A3(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(new_n298_), .A3(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G127gat), .B(G134gat), .Z(new_n306_));
  XOR2_X1   g105(.A(G113gat), .B(G120gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n304_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n297_), .A2(new_n298_), .A3(new_n302_), .A4(new_n310_), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n305_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n309_), .B1(new_n305_), .B2(new_n311_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n272_), .B(new_n282_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT81), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n323_));
  AND2_X1   g122(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n321_), .B(new_n322_), .C1(new_n323_), .C2(new_n324_), .ZN(new_n325_));
  AND3_X1   g124(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n326_));
  INV_X1    g125(.A(G141gat), .ZN(new_n327_));
  INV_X1    g126(.A(G148gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(KEYINPUT3), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(G141gat), .B2(G148gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n326_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT84), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n325_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n325_), .B2(new_n332_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n318_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n315_), .A2(KEYINPUT1), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n317_), .B1(new_n316_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n321_), .A2(new_n322_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n327_), .A2(new_n328_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n336_), .A2(new_n337_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT28), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n336_), .A2(new_n346_), .A3(new_n349_), .A4(new_n337_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G22gat), .B(G50gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n352_), .B(KEYINPUT85), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT89), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n348_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT90), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n348_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n353_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT89), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(G233gat), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT87), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n366_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT88), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n337_), .B1(new_n336_), .B2(new_n346_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n372_), .A2(new_n214_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n367_), .A2(KEYINPUT88), .A3(new_n368_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n371_), .B(new_n374_), .C1(new_n372_), .C2(new_n214_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT90), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n355_), .A2(new_n356_), .A3(new_n379_), .A4(new_n357_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n359_), .A2(new_n362_), .A3(new_n378_), .A4(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n362_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n360_), .A2(new_n361_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n379_), .B1(new_n383_), .B2(new_n356_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n380_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n314_), .B1(new_n381_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n318_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n325_), .A2(new_n332_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT84), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n325_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n388_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n344_), .A2(new_n345_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n309_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n336_), .A2(new_n346_), .A3(new_n308_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(KEYINPUT4), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n398_), .B(new_n309_), .C1(new_n392_), .C2(new_n394_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT92), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n308_), .B1(new_n336_), .B2(new_n346_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(KEYINPUT92), .A3(new_n398_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n397_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G1gat), .B(G29gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT93), .B(G85gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n410_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT95), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n408_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n415_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n417_), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n422_));
  AOI211_X1 g221(.A(new_n415_), .B(new_n408_), .C1(new_n404_), .C2(new_n406_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n424_), .A3(KEYINPUT96), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n422_), .A2(new_n423_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n410_), .A2(new_n417_), .A3(new_n415_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n387_), .A2(new_n425_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n386_), .A2(new_n381_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n273_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n276_), .A2(new_n280_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n432_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n427_), .A2(new_n428_), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n410_), .A2(KEYINPUT33), .A3(new_n415_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n251_), .A2(new_n254_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n247_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n213_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n226_), .A2(new_n232_), .B1(new_n236_), .B2(new_n242_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n277_), .B1(new_n441_), .B2(new_n214_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n258_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n269_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n275_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n273_), .A2(new_n264_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n395_), .A2(new_n396_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n451_), .A2(KEYINPUT94), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n406_), .B1(new_n451_), .B2(KEYINPUT94), .ZN(new_n453_));
  OAI221_X1 g252(.A(new_n419_), .B1(new_n404_), .B2(new_n406_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n437_), .A2(new_n448_), .A3(new_n450_), .A4(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n431_), .B1(new_n436_), .B2(new_n456_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n447_), .A2(new_n203_), .B1(new_n274_), .B2(new_n281_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n386_), .A2(new_n458_), .A3(new_n381_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(new_n429_), .A3(new_n425_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n312_), .A2(new_n313_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n430_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT72), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G232gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT34), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT35), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT68), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT68), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n469_), .A3(KEYINPUT35), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT71), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G29gat), .B(G36gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT69), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n476_), .A2(KEYINPUT69), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n475_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(new_n477_), .A3(new_n474_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n482_), .A3(KEYINPUT15), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT15), .B1(new_n480_), .B2(new_n482_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT65), .B(KEYINPUT6), .Z(new_n487_));
  INV_X1    g286(.A(G99gat), .ZN(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT64), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(G92gat), .B1(KEYINPUT9), .B2(G85gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500_));
  INV_X1    g299(.A(G85gat), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT10), .B(G99gat), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n504_), .A2(G106gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n495_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT66), .A4(KEYINPUT7), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n488_), .A2(new_n489_), .B1(KEYINPUT66), .B2(KEYINPUT7), .ZN(new_n509_));
  OR2_X1    g308(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n492_), .A2(new_n494_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G85gat), .B(G92gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT8), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n508_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n494_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n493_), .A2(new_n490_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT8), .ZN(new_n519_));
  INV_X1    g318(.A(new_n513_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n507_), .B1(new_n514_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n473_), .B1(new_n486_), .B2(new_n522_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n512_), .A2(KEYINPUT8), .A3(new_n513_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n519_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n506_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n480_), .A2(new_n482_), .ZN(new_n527_));
  OAI22_X1  g326(.A1(new_n526_), .A2(new_n527_), .B1(KEYINPUT35), .B2(new_n466_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n464_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n466_), .A2(KEYINPUT35), .ZN(new_n530_));
  INV_X1    g329(.A(new_n527_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n522_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n485_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n483_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n526_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n532_), .A2(new_n535_), .A3(KEYINPUT72), .A4(new_n473_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT70), .B1(new_n486_), .B2(new_n522_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(new_n526_), .A3(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n540_), .A3(new_n532_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n471_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT36), .ZN(new_n544_));
  XOR2_X1   g343(.A(G190gat), .B(G218gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(G134gat), .B(G162gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n529_), .A2(new_n536_), .B1(new_n541_), .B2(new_n471_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(KEYINPUT36), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n537_), .A2(KEYINPUT36), .A3(new_n542_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n548_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n463_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G230gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT11), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(KEYINPUT11), .ZN(new_n560_));
  XOR2_X1   g359(.A(G71gat), .B(G78gat), .Z(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n560_), .A2(new_n561_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n526_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n522_), .A2(new_n564_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(KEYINPUT12), .ZN(new_n568_));
  OR3_X1    g367(.A1(new_n522_), .A2(KEYINPUT12), .A3(new_n564_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n557_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n567_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n570_), .B1(new_n557_), .B2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G120gat), .B(G148gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n572_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n556_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n570_), .B2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(new_n579_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n579_), .B1(new_n578_), .B2(new_n582_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G15gat), .B(G22gat), .ZN(new_n587_));
  INV_X1    g386(.A(G8gat), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G1gat), .B(G8gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(new_n564_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  OR3_X1    g401(.A1(new_n596_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(KEYINPUT17), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n596_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT75), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n531_), .A2(new_n592_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n592_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(new_n527_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G113gat), .B(G141gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G169gat), .B(G197gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n615_), .B(new_n616_), .Z(new_n617_));
  NOR2_X1   g416(.A1(new_n486_), .A2(new_n592_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n531_), .A2(new_n592_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n609_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n614_), .B(new_n617_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT74), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n608_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n614_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n617_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n621_), .A2(new_n622_), .A3(new_n608_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .A4(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n626_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n627_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n623_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n586_), .A2(new_n607_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n555_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT97), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n429_), .A2(new_n425_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n202_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT76), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n632_), .B(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n463_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n586_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n553_), .A2(KEYINPUT37), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n548_), .B(new_n645_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n643_), .A2(new_n648_), .A3(new_n606_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n642_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n638_), .A2(new_n202_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n653_));
  OAI22_X1  g452(.A1(new_n650_), .A2(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n653_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n639_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n639_), .B2(new_n656_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1324gat));
  NOR3_X1   g459(.A1(new_n650_), .A2(G8gat), .A3(new_n458_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n635_), .B2(new_n458_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n458_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n555_), .A2(KEYINPUT100), .A3(new_n664_), .A4(new_n634_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(G8gat), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT39), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n663_), .A2(new_n668_), .A3(G8gat), .A4(new_n665_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n661_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n670_), .B(new_n672_), .ZN(G1325gat));
  OR3_X1    g472(.A1(new_n650_), .A2(G15gat), .A3(new_n462_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G15gat), .B1(new_n636_), .B2(new_n462_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n676_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(G1326gat));
  INV_X1    g478(.A(G22gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n431_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n637_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n683_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n681_), .A2(new_n680_), .ZN(new_n686_));
  OAI22_X1  g485(.A1(new_n684_), .A2(new_n685_), .B1(new_n650_), .B2(new_n686_), .ZN(G1327gat));
  NOR3_X1   g486(.A1(new_n643_), .A2(new_n553_), .A3(new_n607_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n642_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n638_), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n692_));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n463_), .B2(new_n647_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  INV_X1    g494(.A(new_n462_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n695_), .B(new_n648_), .C1(new_n697_), .C2(new_n430_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n606_), .B(new_n632_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n693_), .B1(new_n699_), .B2(new_n703_), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT104), .B(new_n702_), .C1(new_n694_), .C2(new_n698_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n692_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n702_), .B1(new_n694_), .B2(new_n698_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT44), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n638_), .A2(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n691_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  NAND2_X1  g511(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(G36gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n458_), .B1(new_n707_), .B2(KEYINPUT44), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n706_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n458_), .B(KEYINPUT106), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n717_), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n689_), .A2(new_n720_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n689_), .B2(new_n723_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n713_), .B(new_n716_), .C1(new_n719_), .C2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n692_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n459_), .A2(new_n429_), .A3(new_n425_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n435_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n421_), .A2(new_n424_), .A3(new_n730_), .ZN(new_n731_));
  AOI22_X1  g530(.A1(new_n731_), .A2(new_n455_), .B1(new_n381_), .B2(new_n386_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n462_), .B1(new_n729_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n430_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n695_), .B1(new_n735_), .B2(new_n648_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n698_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n703_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT104), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n707_), .A2(new_n693_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n728_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n718_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G36gat), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n726_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n743_), .A2(new_n714_), .A3(new_n715_), .A4(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n727_), .A2(new_n745_), .ZN(G1329gat));
  OAI21_X1  g545(.A(new_n287_), .B1(new_n689_), .B2(new_n462_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n462_), .A2(new_n287_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n709_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT47), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n747_), .C1(new_n709_), .C2(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1330gat));
  AOI21_X1  g553(.A(G50gat), .B1(new_n690_), .B2(new_n681_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n681_), .A2(G50gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n710_), .B2(new_n756_), .ZN(G1331gat));
  NAND4_X1  g556(.A1(new_n555_), .A2(new_n607_), .A3(new_n643_), .A4(new_n641_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n638_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G57gat), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n648_), .A2(new_n606_), .A3(new_n586_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT109), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n463_), .A2(new_n632_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n759_), .A2(G57gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n760_), .B1(new_n764_), .B2(new_n765_), .ZN(G1332gat));
  OAI21_X1  g565(.A(G64gat), .B1(new_n758_), .B2(new_n721_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT48), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n721_), .A2(G64gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n764_), .B2(new_n769_), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n758_), .B2(new_n462_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT49), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n462_), .A2(G71gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n764_), .B2(new_n773_), .ZN(G1334gat));
  OAI21_X1  g573(.A(G78gat), .B1(new_n758_), .B2(new_n431_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT50), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n431_), .A2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n764_), .B2(new_n777_), .ZN(G1335gat));
  NOR2_X1   g577(.A1(new_n586_), .A2(new_n607_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(new_n632_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n699_), .A2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT110), .ZN(new_n783_));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n759_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n780_), .A2(new_n553_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n763_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n501_), .A3(new_n638_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n784_), .A2(new_n788_), .ZN(G1336gat));
  OAI21_X1  g588(.A(G92gat), .B1(new_n783_), .B2(new_n721_), .ZN(new_n790_));
  OR3_X1    g589(.A1(new_n786_), .A2(G92gat), .A3(new_n458_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1337gat));
  NOR3_X1   g591(.A1(new_n786_), .A2(new_n462_), .A3(new_n504_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n782_), .A2(new_n696_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G99gat), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n489_), .A3(new_n681_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n699_), .A2(new_n681_), .A3(new_n781_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n568_), .A2(new_n557_), .A3(new_n569_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n570_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n568_), .A2(new_n569_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n806_), .A3(new_n556_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n580_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n804_), .B1(new_n807_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n556_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n568_), .A2(new_n557_), .A3(new_n569_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(KEYINPUT55), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n577_), .B1(new_n570_), .B2(new_n806_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n811_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n609_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n619_), .A2(new_n610_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n818_), .B(new_n626_), .C1(new_n618_), .C2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n621_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n621_), .A2(new_n820_), .A3(KEYINPUT112), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n572_), .A2(new_n577_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT58), .B1(new_n817_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT113), .B1(new_n647_), .B2(new_n826_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n815_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n814_), .B2(new_n815_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n644_), .A4(new_n646_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n817_), .A2(KEYINPUT58), .A3(new_n825_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n827_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n628_), .A2(new_n631_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n829_), .A2(KEYINPUT111), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n816_), .B1(new_n829_), .B2(KEYINPUT111), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n578_), .A2(new_n582_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n823_), .A2(new_n824_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(KEYINPUT57), .A3(new_n553_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  INV_X1    g646(.A(new_n844_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n811_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n838_), .A3(new_n816_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n848_), .B1(new_n851_), .B2(new_n837_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n847_), .B1(new_n852_), .B2(new_n554_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n836_), .A2(new_n846_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n606_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n641_), .A2(new_n586_), .A3(new_n607_), .A4(new_n647_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT54), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n638_), .A2(new_n387_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861_), .B2(new_n632_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(KEYINPUT59), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT114), .B(KEYINPUT59), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n866_), .B(new_n867_), .C1(new_n860_), .C2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n860_), .A2(new_n868_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT115), .B1(new_n870_), .B2(new_n865_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(G113gat), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n641_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n862_), .B1(new_n872_), .B2(new_n874_), .ZN(G1340gat));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n586_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n861_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n876_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n870_), .A2(new_n586_), .A3(new_n865_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n876_), .ZN(G1341gat));
  AOI21_X1  g679(.A(G127gat), .B1(new_n861_), .B2(new_n607_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n607_), .A2(G127gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT116), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n872_), .B2(new_n883_), .ZN(G1342gat));
  AOI21_X1  g683(.A(G134gat), .B1(new_n861_), .B2(new_n554_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT117), .B(G134gat), .Z(new_n886_));
  NOR2_X1   g685(.A1(new_n647_), .A2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n872_), .B2(new_n887_), .ZN(G1343gat));
  NOR2_X1   g687(.A1(new_n431_), .A2(new_n696_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n858_), .A2(new_n889_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n890_), .A2(new_n759_), .A3(new_n722_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n632_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT118), .B(G141gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1344gat));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n643_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g695(.A1(new_n891_), .A2(new_n607_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1346gat));
  INV_X1    g698(.A(new_n891_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G162gat), .B1(new_n900_), .B2(new_n647_), .ZN(new_n901_));
  INV_X1    g700(.A(G162gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n891_), .A2(new_n902_), .A3(new_n554_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1347gat));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  INV_X1    g704(.A(new_n632_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n638_), .A2(new_n721_), .A3(new_n681_), .A4(new_n462_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  AOI211_X1 g707(.A(new_n906_), .B(new_n908_), .C1(new_n855_), .C2(new_n857_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n905_), .B1(new_n909_), .B2(new_n220_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n858_), .A2(new_n907_), .ZN(new_n911_));
  OAI211_X1 g710(.A(KEYINPUT62), .B(G169gat), .C1(new_n911_), .C2(new_n906_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n909_), .A2(new_n237_), .A3(new_n241_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n910_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT119), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n910_), .A2(new_n912_), .A3(new_n913_), .A4(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1348gat));
  NOR3_X1   g717(.A1(new_n911_), .A2(new_n221_), .A3(new_n586_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n919_), .A2(KEYINPUT121), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(KEYINPUT121), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n221_), .B1(new_n911_), .B2(new_n586_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n923_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n920_), .A2(new_n921_), .B1(new_n924_), .B2(new_n925_), .ZN(G1349gat));
  OR3_X1    g725(.A1(new_n911_), .A2(new_n227_), .A3(new_n606_), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n927_), .A2(KEYINPUT122), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n908_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n929_));
  AOI21_X1  g728(.A(G183gat), .B1(new_n929_), .B2(new_n607_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n927_), .A2(KEYINPUT122), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n928_), .B1(new_n930_), .B2(new_n931_), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n929_), .A2(new_n249_), .A3(new_n554_), .ZN(new_n933_));
  INV_X1    g732(.A(G190gat), .ZN(new_n934_));
  AOI211_X1 g733(.A(KEYINPUT123), .B(new_n934_), .C1(new_n929_), .C2(new_n648_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n858_), .A2(new_n648_), .A3(new_n907_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(G190gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n933_), .B1(new_n935_), .B2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT124), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n941_), .B(new_n933_), .C1(new_n935_), .C2(new_n938_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(G1351gat));
  NOR2_X1   g742(.A1(new_n638_), .A2(new_n721_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n890_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n632_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n949_));
  INV_X1    g748(.A(new_n890_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(new_n944_), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n949_), .B(G204gat), .C1(new_n951_), .C2(new_n586_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n890_), .A2(new_n586_), .A3(new_n945_), .ZN(new_n953_));
  INV_X1    g752(.A(G204gat), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT125), .B1(new_n953_), .B2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n952_), .A2(new_n955_), .ZN(new_n956_));
  NAND4_X1  g755(.A1(new_n950_), .A2(new_n954_), .A3(new_n643_), .A4(new_n944_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n953_), .A2(KEYINPUT126), .A3(new_n954_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n956_), .A2(new_n961_), .ZN(G1353gat));
  AOI211_X1 g761(.A(KEYINPUT63), .B(G211gat), .C1(new_n946_), .C2(new_n607_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n951_), .A2(new_n606_), .ZN(new_n964_));
  XOR2_X1   g763(.A(KEYINPUT63), .B(G211gat), .Z(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n964_), .B2(new_n965_), .ZN(G1354gat));
  NAND2_X1  g765(.A1(new_n946_), .A2(new_n554_), .ZN(new_n967_));
  XOR2_X1   g766(.A(KEYINPUT127), .B(G218gat), .Z(new_n968_));
  NOR2_X1   g767(.A1(new_n647_), .A2(new_n968_), .ZN(new_n969_));
  AOI22_X1  g768(.A1(new_n967_), .A2(new_n968_), .B1(new_n946_), .B2(new_n969_), .ZN(G1355gat));
endmodule


