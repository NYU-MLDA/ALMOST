//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(G141gat), .ZN(new_n205_));
  INV_X1    g004(.A(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT86), .ZN(new_n208_));
  OR3_X1    g007(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT3), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT87), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT2), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n207_), .B1(new_n208_), .B2(KEYINPUT3), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n211_), .A2(KEYINPUT2), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n203_), .B(new_n204_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n203_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT85), .B1(new_n203_), .B2(KEYINPUT1), .ZN(new_n218_));
  OAI221_X1 g017(.A(new_n204_), .B1(KEYINPUT1), .B2(new_n203_), .C1(new_n217_), .C2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(new_n207_), .A3(new_n210_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n202_), .B1(new_n221_), .B2(KEYINPUT29), .ZN(new_n222_));
  INV_X1    g021(.A(G204gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT90), .B1(new_n223_), .B2(G197gat), .ZN(new_n224_));
  INV_X1    g023(.A(G197gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(G204gat), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n223_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT21), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT91), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n230_), .B1(G197gat), .B2(new_n223_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n225_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n231_), .A2(new_n232_), .B1(G197gat), .B2(new_n223_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n228_), .B(new_n229_), .C1(new_n233_), .C2(KEYINPUT21), .ZN(new_n234_));
  INV_X1    g033(.A(new_n229_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(KEYINPUT21), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n222_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT88), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n222_), .A2(new_n240_), .A3(new_n237_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G78gat), .B(G106gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT92), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n242_), .A2(KEYINPUT92), .A3(new_n243_), .A4(new_n245_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G22gat), .B(G50gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT28), .B1(new_n221_), .B2(KEYINPUT29), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n221_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n253_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n254_), .A3(new_n252_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n251_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n250_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT93), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n250_), .A2(new_n261_), .A3(KEYINPUT93), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT25), .B(G183gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G190gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(G169gat), .B2(G176gat), .ZN(new_n271_));
  INV_X1    g070(.A(G169gat), .ZN(new_n272_));
  INV_X1    g071(.A(G176gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n268_), .A2(new_n269_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n276_));
  INV_X1    g075(.A(G183gat), .ZN(new_n277_));
  INV_X1    g076(.A(G190gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT23), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT83), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(G183gat), .A3(G190gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n275_), .B(new_n276_), .C1(new_n280_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n282_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(G183gat), .B2(G190gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(G169gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n267_), .B1(new_n290_), .B2(new_n237_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n276_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT94), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n275_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n280_), .A2(new_n283_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n288_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n291_), .B1(new_n299_), .B2(new_n237_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G226gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT19), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n290_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n237_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n267_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n298_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT95), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n295_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n294_), .A2(KEYINPUT95), .A3(new_n275_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n307_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n306_), .B1(new_n311_), .B2(new_n305_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n303_), .B1(new_n312_), .B2(new_n302_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G8gat), .B(G36gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT18), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(KEYINPUT32), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n311_), .A2(new_n305_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n302_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n291_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(KEYINPUT32), .ZN(new_n322_));
  INV_X1    g121(.A(new_n312_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n321_), .B(new_n322_), .C1(new_n323_), .C2(new_n320_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT96), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327_));
  XOR2_X1   g126(.A(G127gat), .B(G134gat), .Z(new_n328_));
  XOR2_X1   g127(.A(G113gat), .B(G120gat), .Z(new_n329_));
  OR2_X1    g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT84), .B1(new_n328_), .B2(new_n329_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n221_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n328_), .B(new_n329_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n216_), .A2(new_n220_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n327_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT4), .B1(new_n221_), .B2(new_n332_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n326_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n335_), .A3(new_n325_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G1gat), .B(G29gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G57gat), .B(G85gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  NAND3_X1  g143(.A1(new_n338_), .A2(new_n339_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n318_), .B(new_n324_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n321_), .B1(new_n323_), .B2(new_n320_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n317_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n317_), .B(new_n321_), .C1(new_n323_), .C2(new_n320_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT33), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n345_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n326_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n333_), .A2(new_n335_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(KEYINPUT98), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(KEYINPUT98), .B2(new_n357_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n344_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n325_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n338_), .A2(new_n339_), .A3(KEYINPUT33), .A4(new_n344_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n355_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n348_), .B1(new_n353_), .B2(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n247_), .A2(new_n249_), .A3(new_n259_), .A4(new_n257_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n266_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n250_), .A2(new_n261_), .A3(KEYINPUT93), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT93), .B1(new_n250_), .B2(new_n261_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n366_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n346_), .A2(new_n347_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n313_), .A2(new_n350_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n352_), .A2(new_n373_), .A3(KEYINPUT27), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT99), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT99), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n352_), .A2(new_n373_), .A3(new_n376_), .A4(KEYINPUT27), .ZN(new_n377_));
  INV_X1    g176(.A(new_n353_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n375_), .B(new_n377_), .C1(new_n378_), .C2(KEYINPUT27), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n367_), .B1(new_n372_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n381_), .B(G43gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n290_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(new_n332_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(G15gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT30), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT31), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n384_), .A2(new_n389_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n380_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n371_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n379_), .A2(new_n397_), .A3(new_n370_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G15gat), .B(G22gat), .ZN(new_n401_));
  INV_X1    g200(.A(G1gat), .ZN(new_n402_));
  INV_X1    g201(.A(G8gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT14), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G1gat), .B(G8gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G29gat), .B(G36gat), .Z(new_n409_));
  XOR2_X1   g208(.A(G43gat), .B(G50gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n411_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n407_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G229gat), .A2(G233gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT81), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT15), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n411_), .B(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(new_n408_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT82), .ZN(new_n423_));
  INV_X1    g222(.A(new_n412_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(new_n417_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n419_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G113gat), .B(G141gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G169gat), .B(G197gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  XNOR2_X1  g228(.A(new_n426_), .B(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n400_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G183gat), .B(G211gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT80), .ZN(new_n433_));
  XOR2_X1   g232(.A(G127gat), .B(G155gat), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT17), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(KEYINPUT17), .B2(new_n438_), .ZN(new_n441_));
  INV_X1    g240(.A(G64gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G57gat), .ZN(new_n443_));
  INV_X1    g242(.A(G57gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G64gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT69), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT11), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n444_), .A2(G64gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n442_), .A2(G57gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT69), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT11), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G71gat), .B(G78gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n449_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  OAI211_X1 g257(.A(KEYINPUT11), .B(new_n456_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(new_n407_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G231gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n441_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n463_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n440_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G85gat), .ZN(new_n469_));
  INV_X1    g268(.A(G92gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n472_), .B(new_n474_), .C1(KEYINPUT65), .C2(KEYINPUT9), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n471_), .A2(KEYINPUT65), .A3(KEYINPUT9), .A4(new_n473_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT6), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n483_));
  INV_X1    g282(.A(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT64), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n487_), .ZN(new_n489_));
  AND4_X1   g288(.A1(new_n475_), .A2(new_n482_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n471_), .A2(new_n473_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n479_), .B1(G99gat), .B2(G106gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n477_), .A2(KEYINPUT6), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n497_));
  NOR2_X1   g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  OAI22_X1  g297(.A1(new_n495_), .A2(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n500_));
  INV_X1    g299(.A(G99gat), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n501_), .B(new_n484_), .C1(new_n497_), .C2(KEYINPUT66), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT66), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n503_), .A2(KEYINPUT7), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n500_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(KEYINPUT66), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(KEYINPUT7), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(KEYINPUT67), .A4(new_n498_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n499_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n494_), .B1(new_n509_), .B2(new_n492_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n508_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n498_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(KEYINPUT7), .A2(new_n512_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n492_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n494_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n490_), .B1(new_n510_), .B2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(new_n421_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT75), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n411_), .B2(new_n518_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT75), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n519_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT76), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n525_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n521_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n482_), .A2(new_n488_), .A3(new_n475_), .A4(new_n489_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n516_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n533_));
  AOI211_X1 g332(.A(new_n492_), .B(new_n494_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n527_), .B1(new_n413_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n520_), .A2(KEYINPUT76), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(new_n525_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G134gat), .B(G162gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(G190gat), .B(G218gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT78), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n542_), .B(KEYINPUT36), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n531_), .A2(new_n538_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT37), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n552_), .A3(new_n549_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n468_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n458_), .A2(KEYINPUT70), .A3(new_n459_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n555_), .A2(KEYINPUT12), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n460_), .A2(new_n439_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n556_), .A2(new_n535_), .A3(new_n557_), .A4(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n518_), .B2(new_n460_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(KEYINPUT12), .A3(new_n555_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT71), .B1(new_n563_), .B2(new_n518_), .ZN(new_n564_));
  AND2_X1   g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n518_), .B2(new_n460_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n562_), .A2(KEYINPUT72), .A3(new_n564_), .A4(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n564_), .A2(new_n561_), .A3(new_n559_), .A4(new_n566_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n518_), .A2(new_n460_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n518_), .A2(new_n460_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n565_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n567_), .A2(new_n570_), .A3(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G120gat), .B(G148gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n575_), .A2(new_n580_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(KEYINPUT13), .A3(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n554_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT100), .B1(new_n431_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n589_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n591_), .A2(new_n400_), .A3(new_n592_), .A4(new_n430_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n402_), .A3(new_n395_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT38), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT102), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n546_), .A2(new_n599_), .A3(new_n549_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n394_), .B2(new_n399_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n588_), .A2(new_n604_), .A3(new_n430_), .A4(new_n467_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n588_), .A2(new_n430_), .A3(new_n467_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT101), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n609_), .A2(new_n395_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n597_), .B(new_n598_), .C1(new_n402_), .C2(new_n610_), .ZN(G1324gat));
  NAND4_X1  g410(.A1(new_n590_), .A2(new_n403_), .A3(new_n379_), .A4(new_n593_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n603_), .A2(new_n379_), .A3(new_n608_), .A4(new_n605_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n613_), .A2(new_n614_), .A3(G8gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n613_), .B2(G8gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT40), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT40), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n612_), .B(new_n620_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n618_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1325gat));
  NAND2_X1  g423(.A1(new_n609_), .A2(new_n392_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G15gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT105), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n628_), .A3(G15gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n629_), .A3(KEYINPUT41), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT41), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n625_), .B2(G15gat), .ZN(new_n632_));
  AOI211_X1 g431(.A(KEYINPUT105), .B(new_n386_), .C1(new_n609_), .C2(new_n392_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n631_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n594_), .A2(new_n386_), .A3(new_n392_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n634_), .A3(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n370_), .B(KEYINPUT106), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n594_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n606_), .A2(new_n608_), .A3(new_n639_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(new_n642_), .A3(G22gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n641_), .B2(G22gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n600_), .A2(new_n601_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n467_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n588_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n431_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n395_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n551_), .A2(new_n553_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n400_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n398_), .B1(new_n380_), .B2(new_n393_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n656_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n660_));
  OAI22_X1  g459(.A1(new_n658_), .A2(new_n654_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n588_), .A2(new_n430_), .A3(new_n468_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n653_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  AOI211_X1 g465(.A(new_n666_), .B(new_n663_), .C1(new_n657_), .C2(new_n661_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n395_), .A2(G29gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n652_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n651_), .A2(new_n671_), .A3(new_n379_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT45), .ZN(new_n673_));
  INV_X1    g472(.A(new_n379_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n665_), .A2(new_n667_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n675_), .B2(new_n671_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  OAI221_X1 g478(.A(new_n673_), .B1(new_n677_), .B2(KEYINPUT46), .C1(new_n675_), .C2(new_n671_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  AND2_X1   g480(.A1(new_n392_), .A2(G43gat), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n668_), .A2(new_n682_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n431_), .A2(new_n650_), .A3(new_n393_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(G43gat), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(KEYINPUT111), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n684_), .A2(new_n687_), .A3(G43gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT47), .B1(new_n683_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n668_), .A2(new_n682_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n691_), .B(new_n692_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1330gat));
  INV_X1    g493(.A(G50gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n651_), .A2(new_n695_), .A3(new_n639_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT112), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n668_), .A2(new_n697_), .A3(new_n370_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G50gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n668_), .B2(new_n370_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(G1331gat));
  NOR2_X1   g500(.A1(new_n658_), .A2(new_n430_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(new_n587_), .A3(new_n554_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(new_n444_), .A3(new_n395_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n400_), .A2(new_n648_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n430_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n587_), .A2(new_n706_), .A3(new_n467_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n705_), .A2(new_n371_), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n708_), .B2(new_n444_), .ZN(G1332gat));
  NOR2_X1   g508(.A1(new_n705_), .A2(new_n707_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n442_), .B1(new_n710_), .B2(new_n379_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n703_), .A2(new_n442_), .A3(new_n379_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1333gat));
  INV_X1    g514(.A(G71gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n710_), .B2(new_n392_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT49), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n703_), .A2(new_n716_), .A3(new_n392_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1334gat));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n710_), .B2(new_n639_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT50), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n703_), .A2(new_n721_), .A3(new_n639_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1335gat));
  NAND3_X1  g524(.A1(new_n702_), .A2(new_n587_), .A3(new_n649_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n469_), .B1(new_n726_), .B2(new_n371_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n587_), .A2(new_n706_), .A3(new_n468_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n657_), .B2(new_n661_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n371_), .A2(new_n469_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT114), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n730_), .B2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT115), .Z(G1336gat));
  OAI21_X1  g533(.A(G92gat), .B1(new_n730_), .B2(new_n674_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n726_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n470_), .A3(new_n379_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1337gat));
  AOI21_X1  g537(.A(new_n501_), .B1(new_n729_), .B2(new_n392_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n739_), .A2(KEYINPUT116), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(KEYINPUT116), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n392_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n736_), .B2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n741_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT51), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n740_), .A2(new_n747_), .A3(new_n741_), .A4(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1338gat));
  NAND3_X1  g548(.A1(new_n736_), .A2(new_n484_), .A3(new_n370_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n729_), .A2(new_n370_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G106gat), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT52), .B(new_n484_), .C1(new_n729_), .C2(new_n370_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT53), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n750_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1339gat));
  NAND3_X1  g558(.A1(new_n554_), .A2(new_n706_), .A3(new_n588_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(KEYINPUT118), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n554_), .A2(new_n588_), .A3(new_n706_), .A4(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n424_), .A2(new_n416_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n417_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(new_n429_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n423_), .A2(new_n767_), .B1(KEYINPUT120), .B2(new_n769_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n769_), .A2(KEYINPUT120), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n426_), .A2(new_n429_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n581_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n567_), .A2(new_n570_), .A3(new_n774_), .ZN(new_n775_));
  AND4_X1   g574(.A1(new_n564_), .A2(new_n561_), .A3(new_n559_), .A4(new_n566_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n564_), .A2(new_n571_), .A3(new_n561_), .A4(new_n559_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(KEYINPUT55), .B1(new_n777_), .B2(new_n565_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n775_), .A2(new_n778_), .A3(KEYINPUT119), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n580_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n775_), .A2(KEYINPUT119), .A3(new_n778_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT119), .B1(new_n775_), .B2(new_n778_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT56), .B(new_n580_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n773_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n654_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT58), .B(new_n773_), .C1(new_n784_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n430_), .A2(new_n581_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n580_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n794_), .B1(new_n797_), .B2(new_n787_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n583_), .A2(new_n772_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n648_), .B(KEYINPUT57), .C1(new_n798_), .C2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n648_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n793_), .A2(new_n800_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n766_), .B1(new_n804_), .B2(new_n468_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n379_), .A2(new_n371_), .A3(new_n393_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n805_), .A2(new_n370_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n805_), .B2(KEYINPUT122), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n370_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n791_), .A2(new_n792_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n467_), .B1(new_n813_), .B2(new_n800_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n812_), .B(new_n806_), .C1(new_n814_), .C2(new_n766_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n814_), .B2(new_n766_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n809_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n811_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n430_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n821_), .B2(new_n820_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n815_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n804_), .A2(new_n468_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n766_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT121), .A3(new_n812_), .A4(new_n806_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(new_n430_), .A3(new_n829_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n819_), .A2(new_n823_), .B1(new_n830_), .B2(new_n820_), .ZN(G1340gat));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n832_));
  AOI21_X1  g631(.A(G120gat), .B1(new_n587_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n832_), .B2(G120gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n825_), .A2(new_n829_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n588_), .B1(new_n811_), .B2(new_n818_), .ZN(new_n836_));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(G1341gat));
  INV_X1    g637(.A(G127gat), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n825_), .A2(new_n829_), .A3(new_n839_), .A4(new_n467_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n468_), .B1(new_n811_), .B2(new_n818_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n839_), .ZN(G1342gat));
  INV_X1    g641(.A(G134gat), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n825_), .A2(new_n829_), .A3(new_n843_), .A4(new_n602_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n654_), .B1(new_n811_), .B2(new_n818_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n843_), .ZN(G1343gat));
  NAND3_X1  g645(.A1(new_n370_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n805_), .A2(new_n379_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n430_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n587_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n467_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1346gat));
  INV_X1    g654(.A(G162gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n848_), .A2(new_n856_), .A3(new_n602_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n848_), .A2(new_n655_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n856_), .ZN(G1347gat));
  NOR2_X1   g658(.A1(new_n674_), .A2(new_n397_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n430_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT124), .Z(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n638_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G169gat), .B1(new_n805_), .B2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT62), .ZN(new_n865_));
  INV_X1    g664(.A(new_n860_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n639_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT125), .B1(new_n805_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n870_), .B(new_n867_), .C1(new_n814_), .C2(new_n766_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT22), .B(G169gat), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n869_), .A2(new_n871_), .A3(new_n430_), .A4(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n865_), .A2(new_n873_), .ZN(G1348gat));
  NAND3_X1  g673(.A1(new_n869_), .A2(new_n871_), .A3(new_n587_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n805_), .A2(new_n370_), .A3(new_n866_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n588_), .A2(new_n273_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n875_), .A2(new_n273_), .B1(new_n876_), .B2(new_n877_), .ZN(G1349gat));
  NOR2_X1   g677(.A1(new_n468_), .A2(new_n268_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n869_), .A2(new_n871_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(new_n467_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n277_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n869_), .A2(new_n871_), .A3(KEYINPUT126), .A4(new_n879_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n882_), .A2(new_n884_), .A3(new_n885_), .ZN(G1350gat));
  NAND4_X1  g685(.A1(new_n869_), .A2(new_n871_), .A3(new_n269_), .A4(new_n602_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n869_), .A2(new_n655_), .A3(new_n871_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n278_), .ZN(G1351gat));
  NOR3_X1   g688(.A1(new_n674_), .A2(new_n372_), .A3(new_n392_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT127), .B1(new_n805_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n893_), .B(new_n890_), .C1(new_n814_), .C2(new_n766_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G197gat), .B1(new_n895_), .B2(new_n430_), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n225_), .B(new_n706_), .C1(new_n892_), .C2(new_n894_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1352gat));
  AND2_X1   g697(.A1(new_n892_), .A2(new_n894_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G204gat), .B1(new_n899_), .B2(new_n588_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n895_), .A2(new_n223_), .A3(new_n587_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1353gat));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n467_), .A2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n895_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n906_), .ZN(new_n908_));
  AOI211_X1 g707(.A(new_n903_), .B(new_n908_), .C1(new_n892_), .C2(new_n894_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1354gat));
  OAI21_X1  g709(.A(G218gat), .B1(new_n899_), .B2(new_n654_), .ZN(new_n911_));
  INV_X1    g710(.A(G218gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n895_), .A2(new_n912_), .A3(new_n602_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1355gat));
endmodule


