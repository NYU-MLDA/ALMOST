//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT8), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G85gat), .B(G92gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT67), .A3(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT7), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n213_), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n212_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n203_), .B1(new_n210_), .B2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n206_), .A2(new_n203_), .A3(new_n209_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT66), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n219_), .B1(new_n226_), .B2(new_n212_), .ZN(new_n227_));
  OR2_X1    g026(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT64), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(KEYINPUT64), .A3(new_n229_), .ZN(new_n232_));
  AOI21_X1  g031(.A(G106gat), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n204_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT9), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT65), .B(G85gat), .Z(new_n236_));
  INV_X1    g035(.A(G92gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(KEYINPUT9), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n225_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n220_), .B2(new_n221_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n235_), .B(new_n239_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  OAI22_X1  g041(.A1(new_n218_), .A2(new_n227_), .B1(new_n233_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G57gat), .B(G64gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n244_), .A2(KEYINPUT11), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(KEYINPUT11), .ZN(new_n246_));
  XOR2_X1   g045(.A(G71gat), .B(G78gat), .Z(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n246_), .A2(new_n247_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n243_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n226_), .A2(new_n212_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n219_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n212_), .A2(new_n222_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n206_), .A2(new_n209_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT8), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n234_), .A2(KEYINPUT9), .B1(new_n236_), .B2(new_n238_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n261_), .A2(new_n226_), .ZN(new_n262_));
  INV_X1    g061(.A(G106gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n232_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n230_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n257_), .A2(new_n260_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n250_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n254_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G230gat), .A2(G233gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT69), .B1(new_n242_), .B2(new_n233_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n265_), .A2(new_n261_), .A3(new_n226_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT68), .B1(new_n218_), .B2(new_n227_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n257_), .A2(new_n260_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(KEYINPUT12), .A3(new_n251_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n268_), .A2(new_n269_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n267_), .A2(new_n252_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(G230gat), .A3(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G120gat), .B(G148gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT5), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G176gat), .B(G204gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n279_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n202_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(KEYINPUT70), .A3(new_n287_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT13), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT13), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT71), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G232gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT34), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G29gat), .B(G36gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n307_), .A2(KEYINPUT74), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G36gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G29gat), .ZN(new_n311_));
  INV_X1    g110(.A(G29gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G36gat), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n311_), .A2(new_n313_), .A3(KEYINPUT74), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G43gat), .B(G50gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n309_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(new_n308_), .B2(new_n314_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n317_), .A2(new_n319_), .A3(KEYINPUT15), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT15), .B1(new_n317_), .B2(new_n319_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n277_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n303_), .A2(new_n304_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n319_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n243_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n324_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n306_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n218_), .A2(new_n227_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n333_), .A2(new_n275_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n322_), .B1(new_n334_), .B2(new_n274_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT73), .B1(new_n335_), .B2(new_n327_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n324_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n305_), .A3(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G190gat), .B(G218gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT75), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G134gat), .B(G162gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT36), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n332_), .A2(new_n338_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT36), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT76), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n330_), .A2(new_n331_), .A3(new_n306_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n305_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT77), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n332_), .A2(new_n338_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n348_), .ZN(new_n355_));
  AOI211_X1 g154(.A(KEYINPUT37), .B(new_n344_), .C1(new_n352_), .C2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n353_), .B2(new_n348_), .ZN(new_n358_));
  AOI211_X1 g157(.A(KEYINPUT77), .B(new_n347_), .C1(new_n332_), .C2(new_n338_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(KEYINPUT78), .A3(new_n355_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n343_), .B(KEYINPUT79), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n332_), .A2(new_n338_), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n356_), .B1(new_n364_), .B2(KEYINPUT37), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G127gat), .B(G155gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT16), .ZN(new_n368_));
  XOR2_X1   g167(.A(G183gat), .B(G211gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT17), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n366_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G15gat), .B(G22gat), .ZN(new_n373_));
  INV_X1    g172(.A(G1gat), .ZN(new_n374_));
  INV_X1    g173(.A(G8gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT14), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G1gat), .B(G8gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n372_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G231gat), .A2(G233gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n380_), .B(new_n381_), .Z(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(new_n251_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n251_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n370_), .A2(new_n371_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n365_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G169gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT84), .B(G190gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(G183gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT23), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n390_), .B1(new_n392_), .B2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT25), .B(G183gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n391_), .A2(KEYINPUT26), .ZN(new_n401_));
  OR2_X1    g200(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G169gat), .ZN(new_n404_));
  INV_X1    g203(.A(G176gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n406_), .A2(KEYINPUT24), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(KEYINPUT24), .A3(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n407_), .A2(new_n409_), .A3(new_n395_), .A4(new_n396_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n398_), .B1(new_n403_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n411_), .B(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G127gat), .B(G134gat), .Z(new_n415_));
  XOR2_X1   g214(.A(G113gat), .B(G120gat), .Z(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n414_), .B(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(G15gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT30), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT31), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n418_), .A2(new_n423_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT92), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT89), .ZN(new_n431_));
  OR2_X1    g230(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G141gat), .A2(G148gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT87), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(KEYINPUT85), .ZN(new_n439_));
  INV_X1    g238(.A(G141gat), .ZN(new_n440_));
  INV_X1    g239(.A(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n440_), .B(new_n441_), .C1(new_n442_), .C2(KEYINPUT3), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n438_), .B(KEYINPUT85), .C1(G141gat), .C2(G148gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n439_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(KEYINPUT88), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n432_), .A2(KEYINPUT87), .A3(new_n433_), .A4(new_n434_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n437_), .A2(new_n445_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G155gat), .A2(G162gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G155gat), .A2(G162gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n454_), .A2(new_n455_), .A3(KEYINPUT1), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n440_), .A2(new_n441_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT1), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n459_), .B(new_n433_), .C1(new_n460_), .C2(new_n453_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n431_), .B1(new_n457_), .B2(new_n463_), .ZN(new_n464_));
  AOI211_X1 g263(.A(KEYINPUT89), .B(new_n462_), .C1(new_n452_), .C2(new_n456_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n430_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT28), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT28), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n468_), .B(new_n430_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G22gat), .B(G50gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n467_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n429_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n457_), .A2(new_n463_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT89), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n462_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n431_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n468_), .B1(new_n479_), .B2(new_n430_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n469_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n470_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n427_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n467_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n474_), .A2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(G228gat), .A2(G233gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n477_), .A2(new_n430_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n488_), .A2(KEYINPUT91), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G197gat), .B(G204gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G211gat), .B(G218gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT21), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n490_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT21), .B1(new_n491_), .B2(KEYINPUT90), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT21), .B(new_n490_), .C1(new_n491_), .C2(KEYINPUT90), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n488_), .B2(KEYINPUT91), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n487_), .B1(new_n489_), .B2(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n496_), .A2(new_n497_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(new_n487_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(new_n479_), .B2(new_n430_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n486_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n474_), .A2(new_n485_), .A3(new_n504_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT26), .B(G190gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n399_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n410_), .A2(new_n511_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n395_), .B(new_n396_), .C1(G183gat), .C2(G190gat), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(KEYINPUT94), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(KEYINPUT94), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n390_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n501_), .A2(new_n512_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n498_), .B2(new_n411_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G226gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT19), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(new_n519_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT95), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT95), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n517_), .A2(new_n519_), .A3(new_n525_), .A4(new_n522_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n521_), .B(KEYINPUT93), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n501_), .B1(new_n512_), .B2(new_n516_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT20), .B1(new_n498_), .B2(new_n411_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G8gat), .B(G36gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT18), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G64gat), .B(G92gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  AND2_X1   g334(.A1(new_n535_), .A2(KEYINPUT32), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n528_), .A2(new_n529_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n517_), .A2(new_n519_), .ZN(new_n539_));
  OAI22_X1  g338(.A1(new_n538_), .A2(new_n527_), .B1(new_n522_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n536_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G1gat), .B(G29gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G85gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(KEYINPUT98), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G225gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n476_), .A2(new_n478_), .A3(new_n417_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT96), .ZN(new_n553_));
  INV_X1    g352(.A(new_n417_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(new_n477_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n476_), .A2(new_n553_), .A3(new_n478_), .A4(new_n417_), .ZN(new_n557_));
  AOI211_X1 g356(.A(new_n549_), .B(new_n551_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n464_), .A2(new_n465_), .A3(new_n554_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT96), .B1(new_n475_), .B2(new_n417_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n557_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT98), .B1(new_n561_), .B2(new_n550_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n464_), .A2(new_n465_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n560_), .B1(new_n564_), .B2(new_n417_), .ZN(new_n565_));
  NOR4_X1   g364(.A1(new_n464_), .A2(new_n465_), .A3(KEYINPUT96), .A4(new_n554_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT4), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n552_), .A2(KEYINPUT4), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n551_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n548_), .B1(new_n563_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n550_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n549_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n561_), .A2(KEYINPUT98), .A3(new_n550_), .ZN(new_n574_));
  AND4_X1   g373(.A1(new_n548_), .A2(new_n570_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n543_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n570_), .A2(new_n573_), .A3(new_n548_), .A4(new_n574_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(KEYINPUT33), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n535_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n531_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n524_), .A2(new_n530_), .A3(new_n535_), .A4(new_n526_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n568_), .B1(new_n561_), .B2(KEYINPUT4), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n548_), .B1(new_n585_), .B2(new_n550_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n557_), .B(KEYINPUT100), .C1(new_n559_), .C2(new_n560_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT100), .B1(new_n556_), .B2(new_n557_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n551_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n584_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n579_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n563_), .A2(new_n548_), .A3(new_n570_), .A4(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n580_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n508_), .B1(new_n576_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n548_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n573_), .A2(new_n574_), .ZN(new_n597_));
  AOI211_X1 g396(.A(new_n550_), .B(new_n568_), .C1(new_n561_), .C2(KEYINPUT4), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n474_), .A2(new_n485_), .A3(new_n504_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n504_), .B1(new_n474_), .B2(new_n485_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n599_), .B(new_n577_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT27), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n584_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n540_), .A2(new_n581_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(KEYINPUT27), .A3(new_n583_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n426_), .B1(new_n595_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n508_), .B2(new_n607_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n600_), .A2(new_n601_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n604_), .A2(new_n606_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(KEYINPUT101), .A3(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n571_), .A2(new_n575_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n426_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n611_), .A2(new_n614_), .A3(new_n615_), .A4(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n609_), .A2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n388_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n326_), .A2(new_n379_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT81), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n326_), .A2(new_n379_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT82), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n323_), .A2(new_n379_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n621_), .A2(new_n627_), .A3(new_n625_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G113gat), .B(G141gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT83), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G169gat), .B(G197gat), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n631_), .B(new_n632_), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n629_), .B(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n300_), .A2(new_n619_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n615_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n374_), .A3(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT38), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n295_), .A2(new_n634_), .A3(new_n297_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n609_), .B2(new_n617_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n352_), .A2(new_n355_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n344_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n387_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n640_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n615_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n638_), .A2(new_n648_), .ZN(G1324gat));
  OAI21_X1  g448(.A(G8gat), .B1(new_n647_), .B2(new_n613_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(KEYINPUT102), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT39), .B1(new_n650_), .B2(KEYINPUT102), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n635_), .A2(new_n375_), .A3(new_n607_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n653_), .A2(KEYINPUT40), .A3(new_n654_), .A4(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1325gat));
  AOI21_X1  g459(.A(new_n420_), .B1(new_n646_), .B2(new_n616_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n635_), .A2(new_n420_), .A3(new_n616_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1326gat));
  NOR2_X1   g464(.A1(new_n612_), .A2(G22gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT104), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n635_), .A2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G22gat), .B1(new_n647_), .B2(new_n612_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n643_), .A2(new_n386_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n640_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n636_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n639_), .A2(new_n386_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n580_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n542_), .B1(new_n599_), .B2(new_n577_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n612_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n615_), .A2(new_n508_), .A3(new_n613_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n616_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  AND4_X1   g482(.A1(new_n615_), .A2(new_n611_), .A3(new_n616_), .A4(new_n614_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n365_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT43), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n618_), .A2(new_n687_), .A3(new_n365_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n678_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(KEYINPUT44), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n618_), .A2(new_n687_), .A3(new_n365_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n687_), .B1(new_n618_), .B2(new_n365_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n677_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT105), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n691_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT44), .B(new_n677_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n615_), .A2(new_n312_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n676_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n640_), .A2(new_n310_), .A3(new_n607_), .A4(new_n673_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT107), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(KEYINPUT107), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n707_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(KEYINPUT45), .A3(new_n705_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n613_), .B1(new_n689_), .B2(KEYINPUT44), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(new_n691_), .B2(new_n696_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G36gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n711_), .B1(new_n714_), .B2(KEYINPUT106), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n713_), .A2(new_n718_), .A3(G36gat), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .A4(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n698_), .A2(new_n607_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n690_), .B1(new_n689_), .B2(KEYINPUT44), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n694_), .A2(KEYINPUT105), .A3(new_n695_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT106), .B1(new_n724_), .B2(new_n310_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n708_), .A2(new_n710_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n719_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n716_), .A2(new_n717_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n720_), .A2(new_n730_), .ZN(G1329gat));
  NAND3_X1  g530(.A1(new_n700_), .A2(G43gat), .A3(new_n616_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G43gat), .B1(new_n675_), .B2(new_n616_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n732_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1330gat));
  NOR3_X1   g538(.A1(new_n697_), .A2(new_n612_), .A3(new_n699_), .ZN(new_n740_));
  INV_X1    g539(.A(G50gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n508_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT109), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n740_), .A2(new_n741_), .B1(new_n674_), .B2(new_n743_), .ZN(G1331gat));
  INV_X1    g543(.A(new_n634_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n619_), .A2(new_n745_), .A3(new_n298_), .ZN(new_n746_));
  INV_X1    g545(.A(G57gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n636_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n299_), .A2(new_n618_), .A3(new_n745_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(new_n645_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n636_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n751_), .B2(new_n747_), .ZN(G1332gat));
  INV_X1    g551(.A(G64gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n746_), .A2(new_n753_), .A3(new_n607_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n750_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G64gat), .B1(new_n755_), .B2(new_n613_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(KEYINPUT48), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT48), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1333gat));
  INV_X1    g558(.A(G71gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n746_), .A2(new_n760_), .A3(new_n616_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n750_), .A2(new_n616_), .ZN(new_n762_));
  XOR2_X1   g561(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(G71gat), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G71gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(G1334gat));
  INV_X1    g565(.A(G78gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n746_), .A2(new_n767_), .A3(new_n508_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G78gat), .B1(new_n755_), .B2(new_n612_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(G1335gat));
  AND2_X1   g571(.A1(new_n749_), .A2(new_n673_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n636_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n686_), .A2(new_n688_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n298_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n776_), .A2(new_n386_), .A3(new_n634_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT111), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n636_), .A2(new_n236_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT112), .Z(new_n781_));
  AOI21_X1  g580(.A(new_n774_), .B1(new_n779_), .B2(new_n781_), .ZN(G1336gat));
  NAND3_X1  g581(.A1(new_n773_), .A2(new_n237_), .A3(new_n607_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n779_), .A2(new_n607_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n237_), .ZN(G1337gat));
  OAI211_X1 g584(.A(new_n773_), .B(new_n616_), .C1(new_n264_), .C2(new_n230_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT113), .ZN(new_n787_));
  OAI21_X1  g586(.A(G99gat), .B1(new_n778_), .B2(new_n426_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n786_), .B(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n788_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(new_n794_), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n773_), .A2(new_n263_), .A3(new_n508_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n775_), .A2(new_n508_), .A3(new_n777_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G106gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g601(.A1(new_n388_), .A2(new_n745_), .A3(new_n776_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n388_), .A2(new_n745_), .A3(new_n776_), .A4(new_n804_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n278_), .A2(new_n254_), .A3(new_n267_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n269_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n279_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n813_), .B2(KEYINPUT115), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n279_), .B2(new_n812_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n810_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n269_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n279_), .A2(new_n819_), .A3(new_n812_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n814_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n285_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n285_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n634_), .B(new_n287_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n629_), .A2(new_n633_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n633_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n625_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n621_), .A2(new_n627_), .A3(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n827_), .B(new_n829_), .C1(new_n624_), .C2(new_n828_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n826_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n825_), .B1(new_n294_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n831_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(KEYINPUT117), .A3(new_n293_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n824_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n643_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n822_), .A2(new_n823_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n839_), .A2(KEYINPUT58), .A3(new_n287_), .A4(new_n833_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n287_), .B(new_n833_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n843_), .A3(new_n365_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n835_), .A2(KEYINPUT57), .A3(new_n643_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n838_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n387_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n809_), .A2(new_n847_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n611_), .A2(new_n616_), .A3(new_n614_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n849_), .A2(new_n850_), .A3(new_n636_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n844_), .A2(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n840_), .A2(new_n843_), .A3(KEYINPUT118), .A4(new_n365_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n838_), .A3(new_n855_), .A4(new_n845_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n387_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n809_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n858_), .A2(new_n636_), .A3(new_n849_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n634_), .B(new_n852_), .C1(new_n859_), .C2(new_n850_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G113gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n808_), .B1(new_n856_), .B2(new_n387_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n615_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n849_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT119), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n866_), .A3(new_n849_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n745_), .A2(G113gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n861_), .A2(new_n869_), .ZN(G1340gat));
  OAI211_X1 g669(.A(new_n299_), .B(new_n852_), .C1(new_n859_), .C2(new_n850_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G120gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n776_), .A2(KEYINPUT60), .ZN(new_n873_));
  MUX2_X1   g672(.A(new_n873_), .B(KEYINPUT60), .S(G120gat), .Z(new_n874_));
  NAND3_X1  g673(.A1(new_n865_), .A2(new_n867_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(G1341gat));
  OAI211_X1 g675(.A(new_n386_), .B(new_n852_), .C1(new_n859_), .C2(new_n850_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G127gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n387_), .A2(G127gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n865_), .A2(new_n867_), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1342gat));
  NAND3_X1  g680(.A1(new_n865_), .A2(new_n644_), .A3(new_n867_), .ZN(new_n882_));
  INV_X1    g681(.A(G134gat), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n864_), .A2(KEYINPUT59), .B1(new_n848_), .B2(new_n851_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n365_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT120), .B(G134gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n882_), .A2(new_n883_), .B1(new_n884_), .B2(new_n887_), .ZN(G1343gat));
  NOR3_X1   g687(.A1(new_n612_), .A2(new_n607_), .A3(new_n616_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n863_), .A2(new_n634_), .A3(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT121), .B(G141gat), .ZN(new_n891_));
  XOR2_X1   g690(.A(new_n890_), .B(new_n891_), .Z(G1344gat));
  NAND3_X1  g691(.A1(new_n863_), .A2(new_n299_), .A3(new_n889_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT122), .B(G148gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n893_), .B(new_n894_), .Z(G1345gat));
  NAND4_X1  g694(.A1(new_n858_), .A2(new_n636_), .A3(new_n386_), .A4(new_n889_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n863_), .A2(KEYINPUT123), .A3(new_n386_), .A4(new_n889_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n898_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1346gat));
  INV_X1    g702(.A(G162gat), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n863_), .A2(new_n904_), .A3(new_n644_), .A4(new_n889_), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n863_), .A2(new_n365_), .A3(new_n889_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n904_), .ZN(G1347gat));
  AOI21_X1  g706(.A(new_n508_), .B1(new_n809_), .B2(new_n847_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT22), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n613_), .A2(new_n426_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n615_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n908_), .A2(new_n909_), .A3(new_n634_), .A4(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(new_n916_));
  AND4_X1   g715(.A1(new_n634_), .A2(new_n908_), .A3(new_n914_), .A4(new_n912_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n404_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n404_), .B2(new_n916_), .ZN(G1348gat));
  AND2_X1   g718(.A1(new_n908_), .A2(new_n912_), .ZN(new_n920_));
  AOI21_X1  g719(.A(G176gat), .B1(new_n920_), .B2(new_n298_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n862_), .A2(new_n508_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n300_), .A2(new_n405_), .A3(new_n911_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(G1349gat));
  NOR2_X1   g723(.A1(new_n911_), .A2(new_n387_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n908_), .A2(new_n400_), .A3(new_n925_), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT125), .Z(new_n927_));
  AOI21_X1  g726(.A(G183gat), .B1(new_n922_), .B2(new_n925_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1350gat));
  NAND2_X1  g728(.A1(new_n920_), .A2(new_n365_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(G190gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n920_), .A2(new_n644_), .A3(new_n509_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1351gat));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n602_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n858_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n935_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT126), .B1(new_n862_), .B2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT127), .B(G197gat), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n939_), .A2(new_n634_), .A3(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n939_), .B2(new_n634_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1352gat));
  AND2_X1   g742(.A1(new_n936_), .A2(new_n938_), .ZN(new_n944_));
  OAI21_X1  g743(.A(G204gat), .B1(new_n944_), .B2(new_n300_), .ZN(new_n945_));
  INV_X1    g744(.A(G204gat), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n939_), .A2(new_n946_), .A3(new_n299_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1353gat));
  OR2_X1    g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n949_), .B1(new_n939_), .B2(new_n386_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n944_), .A2(new_n387_), .ZN(new_n951_));
  XOR2_X1   g750(.A(KEYINPUT63), .B(G211gat), .Z(new_n952_));
  AOI21_X1  g751(.A(new_n950_), .B1(new_n951_), .B2(new_n952_), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n944_), .B2(new_n885_), .ZN(new_n954_));
  INV_X1    g753(.A(G218gat), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n939_), .A2(new_n955_), .A3(new_n644_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n956_), .ZN(G1355gat));
endmodule


