//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  XOR2_X1   g000(.A(G127gat), .B(G155gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G183gat), .B(G211gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT17), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n208_));
  INV_X1    g007(.A(G231gat), .ZN(new_n209_));
  INV_X1    g008(.A(G233gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n208_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G57gat), .B(G64gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n215_), .B(KEYINPUT11), .Z(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G71gat), .Z(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(G78gat), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n215_), .A2(KEYINPUT11), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n212_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n223_));
  OR3_X1    g022(.A1(new_n214_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225_));
  INV_X1    g024(.A(G1gat), .ZN(new_n226_));
  INV_X1    g025(.A(G8gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT14), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G1gat), .B(G8gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n229_), .B(new_n230_), .Z(new_n231_));
  XOR2_X1   g030(.A(new_n231_), .B(KEYINPUT75), .Z(new_n232_));
  OAI21_X1  g031(.A(new_n222_), .B1(new_n214_), .B2(new_n223_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n224_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n206_), .A2(KEYINPUT17), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n232_), .B1(new_n224_), .B2(new_n233_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT78), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n237_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n235_), .A4(new_n234_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G29gat), .B(G36gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT73), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT73), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n244_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n246_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT15), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT15), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G99gat), .A2(G106gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT6), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(KEYINPUT64), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n263_));
  INV_X1    g062(.A(G99gat), .ZN(new_n264_));
  INV_X1    g063(.A(G106gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n268_));
  OAI22_X1  g067(.A1(new_n266_), .A2(new_n267_), .B1(new_n268_), .B2(new_n260_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n262_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G85gat), .B(G92gat), .Z(new_n271_));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT8), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n272_), .A2(KEYINPUT8), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n270_), .B(new_n274_), .C1(new_n272_), .C2(KEYINPUT8), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT10), .B(G99gat), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n265_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n271_), .A2(KEYINPUT9), .ZN(new_n283_));
  INV_X1    g082(.A(G85gat), .ZN(new_n284_));
  INV_X1    g083(.A(G92gat), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n284_), .A2(new_n285_), .A3(KEYINPUT9), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n282_), .A2(new_n283_), .A3(new_n259_), .A4(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT70), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n280_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n278_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n257_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n277_), .A2(new_n279_), .A3(new_n287_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT35), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G232gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT34), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n292_), .A2(new_n253_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n296_), .A2(new_n293_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT36), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G190gat), .B(G218gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT74), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G134gat), .B(G162gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n299_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n291_), .A2(new_n306_), .A3(new_n297_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n300_), .A2(new_n301_), .A3(new_n305_), .A4(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n305_), .B(KEYINPUT36), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n291_), .A2(new_n306_), .A3(new_n297_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n306_), .B1(new_n291_), .B2(new_n297_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT37), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT37), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n308_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n243_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT79), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G197gat), .B(G204gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT21), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323_));
  INV_X1    g122(.A(G197gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G204gat), .ZN(new_n325_));
  INV_X1    g124(.A(G204gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G197gat), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n325_), .A2(new_n327_), .A3(KEYINPUT94), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT21), .B1(new_n325_), .B2(KEYINPUT94), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n322_), .B(new_n323_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n320_), .A2(new_n321_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(G169gat), .B2(G176gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT85), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(G169gat), .B2(G176gat), .ZN(new_n338_));
  INV_X1    g137(.A(G169gat), .ZN(new_n339_));
  INV_X1    g138(.A(G176gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(KEYINPUT85), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n336_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G183gat), .ZN(new_n344_));
  INV_X1    g143(.A(G183gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT25), .ZN(new_n346_));
  INV_X1    g145(.A(G190gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT26), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT26), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G190gat), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n344_), .A2(new_n346_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n335_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n342_), .A2(new_n351_), .A3(new_n355_), .A4(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G169gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n362_), .B(new_n352_), .C1(G183gat), .C2(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n357_), .A2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT20), .B1(new_n334_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT84), .B1(new_n345_), .B2(KEYINPUT25), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(new_n343_), .A3(G183gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n343_), .B2(G183gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n345_), .A2(KEYINPUT83), .A3(KEYINPUT25), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n367_), .B(new_n342_), .C1(new_n372_), .C2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT24), .B1(new_n341_), .B2(new_n338_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n362_), .A2(new_n352_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT87), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n341_), .A2(new_n338_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n381_), .B(new_n355_), .C1(new_n382_), .C2(KEYINPUT24), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n377_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n348_), .A2(new_n350_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n385_), .A2(new_n371_), .A3(new_n375_), .A4(new_n374_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n367_), .B1(new_n386_), .B2(new_n342_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n364_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n366_), .B1(new_n388_), .B2(new_n334_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n334_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n395_), .B(new_n364_), .C1(new_n384_), .C2(new_n387_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n334_), .B2(new_n365_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n398_), .A3(new_n393_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G8gat), .B(G36gat), .Z(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT18), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n389_), .A2(new_n393_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n396_), .A2(new_n398_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n392_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n409_), .A3(new_n404_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n406_), .A2(KEYINPUT103), .A3(KEYINPUT27), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT103), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(KEYINPUT27), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n404_), .B1(new_n394_), .B2(new_n399_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417_));
  INV_X1    g216(.A(G141gat), .ZN(new_n418_));
  INV_X1    g217(.A(G148gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G141gat), .A2(G148gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT2), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G155gat), .B(G162gat), .Z(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n418_), .A2(new_n419_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n421_), .ZN(new_n431_));
  OR2_X1    g230(.A1(G155gat), .A2(G162gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT1), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n428_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n395_), .B1(KEYINPUT29), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G228gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT93), .ZN(new_n443_));
  OR3_X1    g242(.A1(new_n437_), .A2(new_n443_), .A3(KEYINPUT29), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n437_), .B2(KEYINPUT29), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G22gat), .B(G50gat), .Z(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G78gat), .B(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT95), .ZN(new_n450_));
  INV_X1    g249(.A(new_n447_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n444_), .A2(new_n451_), .A3(new_n445_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n449_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n441_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n456_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n440_), .A3(new_n453_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  AOI211_X1 g259(.A(new_n392_), .B(new_n366_), .C1(new_n388_), .C2(new_n334_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n393_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n405_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n410_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT27), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT104), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n464_), .A2(KEYINPUT104), .A3(new_n465_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n416_), .B(new_n460_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G71gat), .B(G99gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT89), .B(G43gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT88), .B(KEYINPUT30), .Z(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G227gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(G15gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n388_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT91), .ZN(new_n478_));
  INV_X1    g277(.A(new_n476_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n364_), .B(new_n479_), .C1(new_n384_), .C2(new_n387_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n477_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n478_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n473_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT91), .ZN(new_n485_));
  INV_X1    g284(.A(new_n473_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n477_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT31), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n483_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n491_));
  INV_X1    g290(.A(G134gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G127gat), .ZN(new_n493_));
  INV_X1    g292(.A(G127gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G134gat), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n493_), .A2(new_n495_), .A3(KEYINPUT90), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT90), .B1(new_n493_), .B2(new_n495_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G113gat), .B(G120gat), .Z(new_n498_));
  NOR3_X1   g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G120gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n495_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n493_), .A2(new_n495_), .A3(KEYINPUT90), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n500_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OAI22_X1  g304(.A1(new_n490_), .A2(new_n491_), .B1(new_n499_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n483_), .A2(new_n488_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT31), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n499_), .A2(new_n505_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n483_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G1gat), .B(G29gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G57gat), .B(G85gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n427_), .A2(new_n426_), .B1(new_n431_), .B2(new_n435_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n499_), .B2(new_n505_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n503_), .A2(new_n504_), .A3(new_n500_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n498_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n432_), .A2(new_n434_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n425_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n424_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n522_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n429_), .A2(new_n430_), .A3(new_n421_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n427_), .B2(new_n433_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n520_), .B(new_n521_), .C1(new_n529_), .C2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n519_), .A2(new_n532_), .A3(KEYINPUT97), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT97), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n509_), .A2(new_n534_), .A3(new_n437_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G225gat), .A2(G233gat), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT100), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT100), .ZN(new_n539_));
  INV_X1    g338(.A(new_n537_), .ZN(new_n540_));
  AOI211_X1 g339(.A(new_n539_), .B(new_n540_), .C1(new_n533_), .C2(new_n535_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT4), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n509_), .A2(new_n543_), .A3(new_n437_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n537_), .B(KEYINPUT98), .Z(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n517_), .B1(new_n542_), .B2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n540_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT100), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n548_), .A2(new_n517_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n506_), .A2(new_n511_), .A3(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n468_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT101), .B(KEYINPUT33), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n516_), .B1(new_n536_), .B2(new_n546_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n545_), .A2(new_n537_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n560_), .B1(new_n544_), .B2(new_n561_), .ZN(new_n562_));
  OAI211_X1 g361(.A(KEYINPUT33), .B(new_n516_), .C1(new_n544_), .C2(new_n547_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n542_), .B2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n559_), .A2(new_n564_), .A3(new_n464_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n394_), .A2(KEYINPUT32), .A3(new_n404_), .A4(new_n399_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n549_), .A2(new_n553_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n460_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT102), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n554_), .A2(new_n460_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n416_), .B(new_n572_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT102), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n574_), .B(new_n460_), .C1(new_n565_), .C2(new_n569_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n506_), .A2(new_n511_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n557_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n222_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n292_), .A2(KEYINPUT68), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT68), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n277_), .A2(new_n279_), .A3(new_n287_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n581_), .B1(new_n582_), .B2(new_n222_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n580_), .B(new_n583_), .C1(new_n579_), .C2(new_n292_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n222_), .A2(KEYINPUT12), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n292_), .B2(new_n579_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n586_), .B1(new_n292_), .B2(new_n579_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n589_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n587_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G120gat), .B(G148gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G176gat), .B(G204gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n587_), .A2(new_n593_), .A3(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT13), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT13), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n605_), .A3(new_n602_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n252_), .B(KEYINPUT80), .ZN(new_n608_));
  INV_X1    g407(.A(new_n231_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n608_), .A2(new_n609_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n231_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n616_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(G113gat), .B(G141gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT81), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G169gat), .B(G197gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n621_), .B(new_n622_), .Z(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n615_), .A2(new_n619_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n613_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n623_), .B1(new_n626_), .B2(new_n618_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(KEYINPUT82), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT82), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n629_), .B(new_n623_), .C1(new_n626_), .C2(new_n618_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n607_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n578_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n319_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n226_), .A3(new_n554_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n313_), .B(KEYINPUT105), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n578_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n633_), .A2(new_n242_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n555_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n637_), .A2(new_n638_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n639_), .A2(new_n645_), .A3(new_n646_), .ZN(G1324gat));
  OAI21_X1  g446(.A(new_n416_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n635_), .A2(G8gat), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G8gat), .B1(new_n644_), .B2(new_n649_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n654_), .B(new_n655_), .Z(G1325gat));
  INV_X1    g455(.A(new_n577_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n642_), .A2(new_n657_), .A3(new_n643_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(G15gat), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n636_), .A2(new_n475_), .A3(new_n657_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n660_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT108), .Z(G1326gat));
  OAI21_X1  g464(.A(G22gat), .B1(new_n644_), .B2(new_n460_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT42), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n460_), .A2(G22gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n635_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT109), .ZN(G1327gat));
  NOR2_X1   g469(.A1(new_n243_), .A2(new_n313_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n634_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(G29gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n554_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT112), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT113), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT111), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n317_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n314_), .A2(KEYINPUT111), .A3(new_n316_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n578_), .B2(KEYINPUT110), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT110), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n684_), .B(new_n557_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  OR3_X1    g485(.A1(new_n578_), .A2(KEYINPUT43), .A3(new_n317_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n633_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n677_), .A2(KEYINPUT113), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n242_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n678_), .B1(new_n688_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n686_), .A2(new_n687_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n691_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n678_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n693_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n555_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n675_), .B1(new_n697_), .B2(new_n674_), .ZN(G1328gat));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n695_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n691_), .B(new_n678_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n648_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(KEYINPUT114), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n634_), .A2(new_n703_), .A3(new_n648_), .A4(new_n671_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n706_), .A2(KEYINPUT45), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT114), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(KEYINPUT45), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n699_), .B1(new_n705_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n710_), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT46), .B(new_n712_), .C1(new_n702_), .C2(new_n704_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1329gat));
  NAND2_X1  g513(.A1(new_n657_), .A2(G43gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n716_));
  INV_X1    g515(.A(G43gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(new_n672_), .B2(new_n577_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT115), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n716_), .A2(KEYINPUT47), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT47), .B1(new_n716_), .B2(new_n719_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1330gat));
  INV_X1    g521(.A(new_n460_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G50gat), .B1(new_n673_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n692_), .A2(new_n696_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n723_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(G1331gat));
  NAND3_X1  g526(.A1(new_n238_), .A2(new_n631_), .A3(new_n241_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n607_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n642_), .A2(new_n729_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(KEYINPUT116), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(KEYINPUT116), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n554_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n578_), .A2(new_n632_), .A3(new_n607_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n319_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n554_), .A2(new_n734_), .ZN(new_n737_));
  OAI22_X1  g536(.A1(new_n733_), .A2(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(G1332gat));
  OR3_X1    g537(.A1(new_n736_), .A2(G64gat), .A3(new_n649_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n731_), .A2(new_n648_), .A3(new_n732_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(G64gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G64gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT117), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n739_), .B(KEYINPUT117), .C1(new_n742_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1333gat));
  OR3_X1    g547(.A1(new_n736_), .A2(G71gat), .A3(new_n577_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n731_), .A2(new_n657_), .A3(new_n732_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G71gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G71gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1334gat));
  OR3_X1    g553(.A1(new_n736_), .A2(G78gat), .A3(new_n460_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n731_), .A2(new_n723_), .A3(new_n732_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G78gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G78gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n735_), .A2(new_n671_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n284_), .A3(new_n554_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n607_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n242_), .A3(new_n631_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n688_), .A2(new_n555_), .A3(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n763_), .B1(new_n766_), .B2(new_n284_), .ZN(G1336gat));
  NOR3_X1   g566(.A1(new_n688_), .A2(new_n649_), .A3(new_n765_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n648_), .A2(new_n285_), .ZN(new_n769_));
  OAI22_X1  g568(.A1(new_n768_), .A2(new_n285_), .B1(new_n761_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT118), .ZN(G1337gat));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n281_), .A3(new_n657_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n688_), .A2(new_n577_), .A3(new_n765_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(new_n264_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR3_X1   g574(.A1(new_n761_), .A2(G106gat), .A3(new_n460_), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n460_), .B(new_n765_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT52), .B1(new_n777_), .B2(new_n265_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n765_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n693_), .A2(new_n723_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n776_), .B1(new_n778_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n784_), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n776_), .B(new_n786_), .C1(new_n778_), .C2(new_n782_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1339gat));
  INV_X1    g587(.A(new_n317_), .ZN(new_n789_));
  NOR4_X1   g588(.A1(new_n764_), .A2(new_n789_), .A3(KEYINPUT54), .A4(new_n728_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n728_), .B1(new_n606_), .B2(new_n604_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n317_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n790_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n617_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n610_), .A2(new_n795_), .A3(KEYINPUT120), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT120), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n614_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n624_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT121), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n799_), .A2(new_n800_), .A3(KEYINPUT121), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n803_), .A2(new_n625_), .A3(new_n602_), .A4(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n589_), .A2(KEYINPUT55), .A3(new_n591_), .A4(new_n592_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n593_), .A2(new_n807_), .ZN(new_n808_));
  AND4_X1   g607(.A1(new_n583_), .A2(new_n589_), .A3(new_n580_), .A4(new_n591_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n806_), .B(new_n808_), .C1(new_n809_), .C2(new_n585_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n600_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n600_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n805_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT58), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n805_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n600_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n600_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(KEYINPUT122), .A3(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n817_), .A2(new_n789_), .A3(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n628_), .A2(new_n630_), .A3(new_n602_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n603_), .A2(new_n625_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n313_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n825_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n827_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT57), .A3(new_n313_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n824_), .A2(new_n831_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n794_), .B1(new_n836_), .B2(new_n242_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n468_), .A2(new_n555_), .A3(new_n577_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(G113gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n632_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(KEYINPUT123), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n840_), .A2(KEYINPUT123), .A3(KEYINPUT59), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n631_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n842_), .B1(new_n847_), .B2(new_n841_), .ZN(G1340gat));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n607_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT124), .B1(new_n849_), .B2(KEYINPUT60), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n840_), .B(new_n852_), .C1(new_n853_), .C2(new_n850_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n607_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n849_), .ZN(G1341gat));
  NAND3_X1  g655(.A1(new_n840_), .A2(new_n494_), .A3(new_n243_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n242_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n494_), .ZN(G1342gat));
  NAND3_X1  g658(.A1(new_n840_), .A2(new_n492_), .A3(new_n641_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n317_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n492_), .ZN(G1343gat));
  NOR3_X1   g661(.A1(new_n837_), .A2(new_n460_), .A3(new_n657_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n863_), .A2(new_n649_), .A3(new_n554_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(new_n418_), .A3(new_n632_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n649_), .A3(new_n554_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G141gat), .B1(new_n866_), .B2(new_n631_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1344gat));
  NAND3_X1  g667(.A1(new_n864_), .A2(new_n419_), .A3(new_n764_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G148gat), .B1(new_n866_), .B2(new_n607_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1345gat));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  OR3_X1    g671(.A1(new_n866_), .A2(new_n242_), .A3(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n866_), .B2(new_n242_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1346gat));
  NAND2_X1  g674(.A1(new_n864_), .A2(new_n641_), .ZN(new_n876_));
  INV_X1    g675(.A(G162gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n876_), .A2(new_n877_), .B1(new_n864_), .B2(new_n878_), .ZN(G1347gat));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n657_), .A2(new_n460_), .A3(new_n648_), .A4(new_n555_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n631_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n880_), .B1(new_n837_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n834_), .B2(new_n313_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n313_), .ZN(new_n886_));
  AOI211_X1 g685(.A(new_n830_), .B(new_n886_), .C1(new_n833_), .C2(new_n827_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n243_), .B1(new_n888_), .B2(new_n824_), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT125), .B(new_n882_), .C1(new_n889_), .C2(new_n794_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n884_), .A2(new_n890_), .A3(G169gat), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n884_), .A2(new_n890_), .A3(KEYINPUT126), .A4(G169gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(KEYINPUT62), .A3(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n891_), .A2(new_n892_), .A3(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT22), .B(G169gat), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n882_), .B(new_n898_), .C1(new_n889_), .C2(new_n794_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(new_n897_), .A3(new_n899_), .ZN(G1348gat));
  NOR2_X1   g699(.A1(new_n837_), .A2(new_n881_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n764_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G176gat), .ZN(G1349gat));
  NOR3_X1   g702(.A1(new_n837_), .A2(new_n242_), .A3(new_n881_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(G183gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n344_), .A2(new_n346_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n904_), .ZN(G1350gat));
  NAND2_X1  g706(.A1(new_n641_), .A2(new_n385_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT127), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n901_), .A2(new_n909_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n837_), .A2(new_n317_), .A3(new_n881_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n347_), .ZN(G1351gat));
  NOR2_X1   g711(.A1(new_n649_), .A2(new_n554_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n863_), .A2(new_n632_), .A3(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g714(.A1(new_n863_), .A2(new_n764_), .A3(new_n913_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g716(.A(KEYINPUT63), .B(G211gat), .ZN(new_n918_));
  OR2_X1    g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n863_), .A2(new_n243_), .A3(new_n913_), .ZN(new_n920_));
  MUX2_X1   g719(.A(new_n918_), .B(new_n919_), .S(new_n920_), .Z(G1354gat));
  NAND2_X1  g720(.A1(new_n863_), .A2(new_n913_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G218gat), .B1(new_n922_), .B2(new_n317_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n640_), .A2(G218gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(new_n924_), .ZN(G1355gat));
endmodule


