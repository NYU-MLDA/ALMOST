//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G71gat), .B(G78gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n205_));
  INV_X1    g004(.A(new_n203_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT9), .A3(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(KEYINPUT9), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n214_), .A2(new_n218_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n222_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AOI211_X1 g029(.A(KEYINPUT8), .B(new_n226_), .C1(new_n230_), .C2(new_n214_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(G99gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n216_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n212_), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n227_), .B(new_n235_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n226_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n232_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n209_), .B(new_n225_), .C1(new_n231_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT64), .ZN(new_n242_));
  INV_X1    g041(.A(new_n225_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n211_), .A2(new_n213_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n235_), .A2(new_n227_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n239_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT8), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n238_), .A2(new_n232_), .A3(new_n239_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n243_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n209_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n242_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n209_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n225_), .B1(new_n231_), .B2(new_n240_), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n252_), .A2(KEYINPUT65), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(KEYINPUT65), .B2(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G230gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n254_), .B2(new_n253_), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n231_), .A2(new_n240_), .A3(KEYINPUT66), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n225_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n253_), .A2(KEYINPUT12), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n261_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n258_), .B1(new_n249_), .B2(new_n209_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n256_), .A2(new_n258_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT5), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G176gat), .B(G204gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n270_), .B(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n275_), .A2(KEYINPUT13), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT13), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G29gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G43gat), .B(G50gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n249_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G232gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT34), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT66), .B1(new_n231_), .B2(new_n240_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n247_), .A2(new_n263_), .A3(new_n248_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n243_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n281_), .B(KEYINPUT15), .Z(new_n288_));
  OAI221_X1 g087(.A(new_n282_), .B1(KEYINPUT35), .B2(new_n284_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n284_), .A2(KEYINPUT35), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(KEYINPUT68), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n289_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G190gat), .B(G218gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G134gat), .B(G162gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT36), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n295_), .B(KEYINPUT36), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n292_), .A2(new_n299_), .ZN(new_n300_));
  OR3_X1    g099(.A1(new_n297_), .A2(new_n300_), .A3(KEYINPUT37), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n298_), .B(KEYINPUT69), .Z(new_n302_));
  NOR2_X1   g101(.A1(new_n292_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT37), .B1(new_n297_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT17), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G127gat), .B(G155gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT16), .ZN(new_n309_));
  XOR2_X1   g108(.A(G183gat), .B(G211gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n209_), .B(new_n312_), .Z(new_n313_));
  XOR2_X1   g112(.A(G15gat), .B(G22gat), .Z(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT70), .B(G1gat), .Z(new_n315_));
  XOR2_X1   g114(.A(KEYINPUT71), .B(G8gat), .Z(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n314_), .B1(new_n317_), .B2(KEYINPUT14), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G1gat), .B(G8gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n313_), .B(new_n320_), .ZN(new_n321_));
  AOI211_X1 g120(.A(new_n307_), .B(new_n311_), .C1(new_n321_), .C2(KEYINPUT72), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(KEYINPUT72), .B2(new_n321_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n311_), .B(new_n307_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT73), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n321_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n278_), .A2(new_n306_), .A3(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n328_), .B(KEYINPUT74), .Z(new_n329_));
  XOR2_X1   g128(.A(G1gat), .B(G29gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT97), .B(G85gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT0), .B(G57gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  NAND2_X1  g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT83), .ZN(new_n336_));
  XOR2_X1   g135(.A(KEYINPUT84), .B(KEYINPUT2), .Z(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT85), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n341_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(G141gat), .ZN(new_n343_));
  INV_X1    g142(.A(G148gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(KEYINPUT3), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(G141gat), .B2(G148gat), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n340_), .A2(new_n342_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n338_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT86), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G155gat), .ZN(new_n352_));
  INV_X1    g151(.A(G162gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n353_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(KEYINPUT1), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n355_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n360_));
  OAI221_X1 g159(.A(new_n336_), .B1(G141gat), .B2(G148gat), .C1(new_n358_), .C2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G127gat), .B(G134gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G113gat), .B(G120gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n362_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT96), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n362_), .A2(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n362_), .A2(new_n368_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(KEYINPUT4), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n374_), .A2(new_n375_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n372_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n334_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n379_), .A3(new_n334_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT78), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n385_), .A2(KEYINPUT24), .ZN(new_n386_));
  INV_X1    g185(.A(G169gat), .ZN(new_n387_));
  INV_X1    g186(.A(G176gat), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n385_), .B(KEYINPUT24), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT23), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT26), .B(G190gat), .ZN(new_n392_));
  INV_X1    g191(.A(G183gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT25), .B1(new_n393_), .B2(KEYINPUT77), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n393_), .A2(KEYINPUT25), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n392_), .B(new_n394_), .C1(new_n395_), .C2(KEYINPUT77), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n386_), .A2(new_n389_), .A3(new_n391_), .A4(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n391_), .A2(new_n398_), .B1(G169gat), .B2(G176gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT22), .B1(new_n387_), .B2(KEYINPUT79), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n387_), .A2(KEYINPUT22), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n388_), .B(new_n400_), .C1(new_n401_), .C2(KEYINPUT79), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(G15gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT30), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n404_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G71gat), .B(G99gat), .ZN(new_n410_));
  INV_X1    g209(.A(G43gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n409_), .B(new_n412_), .Z(new_n413_));
  XNOR2_X1  g212(.A(new_n368_), .B(KEYINPUT31), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT82), .Z(new_n415_));
  OR2_X1    g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(KEYINPUT82), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n383_), .A2(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n357_), .A2(new_n361_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT29), .ZN(new_n422_));
  XOR2_X1   g221(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n423_), .B1(new_n362_), .B2(KEYINPUT29), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G22gat), .B(G50gat), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n427_), .A2(new_n429_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT88), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n432_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n430_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n362_), .A2(KEYINPUT29), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT21), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G197gat), .B(G204gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT91), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G211gat), .B(G218gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n439_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n438_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n445_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n437_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G228gat), .ZN(new_n448_));
  INV_X1    g247(.A(G233gat), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n449_), .A2(KEYINPUT89), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(KEYINPUT89), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n448_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT90), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n447_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n437_), .A2(new_n453_), .A3(new_n446_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(KEYINPUT92), .Z(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT93), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n455_), .A2(KEYINPUT93), .A3(new_n456_), .A4(new_n458_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n433_), .A2(new_n436_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n434_), .A2(new_n430_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n455_), .A2(new_n456_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n457_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n459_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n464_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n404_), .A2(new_n446_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT25), .B(G183gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n392_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT24), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n384_), .A2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n389_), .A2(new_n391_), .A3(new_n473_), .A4(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT22), .B(G169gat), .Z(new_n477_));
  OAI21_X1  g276(.A(new_n399_), .B1(G176gat), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n471_), .B(KEYINPUT20), .C1(new_n446_), .C2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G226gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT19), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n446_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n484_), .B(KEYINPUT20), .C1(new_n446_), .C2(new_n404_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G8gat), .B(G36gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G64gat), .B(G92gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n492_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n483_), .A2(new_n494_), .A3(new_n486_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT95), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n487_), .A2(KEYINPUT95), .A3(new_n492_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n485_), .A2(new_n482_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n501_), .B1(new_n482_), .B2(new_n480_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n495_), .B(KEYINPUT27), .C1(new_n502_), .C2(new_n494_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n420_), .A2(new_n470_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n383_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n507_), .B(new_n505_), .C1(new_n464_), .C2(new_n469_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n382_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n371_), .A2(new_n372_), .A3(new_n376_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n334_), .B1(new_n378_), .B2(new_n373_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n497_), .A2(new_n498_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n377_), .A2(KEYINPUT33), .A3(new_n379_), .A4(new_n334_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n494_), .A2(KEYINPUT32), .ZN(new_n516_));
  MUX2_X1   g315(.A(new_n502_), .B(new_n487_), .S(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n382_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(new_n380_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n470_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n508_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n506_), .B1(new_n522_), .B2(new_n419_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n320_), .B(new_n281_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n288_), .A2(new_n320_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n320_), .A2(new_n281_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n525_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G169gat), .B(G197gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n527_), .A2(new_n530_), .A3(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n536_), .A2(KEYINPUT75), .A3(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT76), .Z(new_n543_));
  NOR3_X1   g342(.A1(new_n329_), .A2(new_n523_), .A3(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n507_), .A2(new_n315_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n547_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n297_), .A2(new_n300_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n523_), .A2(new_n550_), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n278_), .A2(KEYINPUT100), .A3(new_n542_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n327_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT100), .B1(new_n278_), .B2(new_n542_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(G1gat), .B1(new_n556_), .B2(new_n507_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n548_), .A2(new_n549_), .A3(new_n557_), .ZN(G1324gat));
  INV_X1    g357(.A(new_n316_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n544_), .A2(new_n504_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n504_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT39), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n562_), .A2(new_n563_), .A3(G8gat), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n562_), .B2(G8gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n560_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT40), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT40), .B(new_n560_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(G1325gat));
  INV_X1    g369(.A(new_n419_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n544_), .A2(new_n406_), .A3(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n572_), .B(KEYINPUT101), .Z(new_n573_));
  OAI21_X1  g372(.A(G15gat), .B1(new_n556_), .B2(new_n419_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT41), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(KEYINPUT41), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n573_), .A2(new_n575_), .A3(new_n576_), .ZN(G1326gat));
  INV_X1    g376(.A(G22gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n470_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n544_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n561_), .B2(new_n579_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n580_), .B1(new_n583_), .B2(new_n584_), .ZN(G1327gat));
  NOR2_X1   g384(.A1(new_n523_), .A2(new_n543_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n550_), .A2(new_n327_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n278_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n589_), .A2(G29gat), .A3(new_n507_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT43), .B1(new_n523_), .B2(new_n305_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT43), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n571_), .B1(new_n508_), .B2(new_n521_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n592_), .B(new_n306_), .C1(new_n593_), .C2(new_n506_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n552_), .A2(new_n327_), .A3(new_n554_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT103), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n595_), .A2(KEYINPUT44), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT44), .B1(new_n595_), .B2(new_n598_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT104), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n383_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(G29gat), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n601_), .B2(new_n383_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n590_), .B1(new_n604_), .B2(new_n605_), .ZN(G1328gat));
  INV_X1    g405(.A(G36gat), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n504_), .A2(new_n607_), .ZN(new_n608_));
  OR3_X1    g407(.A1(new_n589_), .A2(KEYINPUT45), .A3(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT45), .B1(new_n589_), .B2(new_n608_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n599_), .A2(new_n600_), .A3(new_n505_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n611_), .B1(new_n612_), .B2(new_n607_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT46), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI211_X1 g414(.A(KEYINPUT46), .B(new_n611_), .C1(new_n612_), .C2(new_n607_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1329gat));
  XNOR2_X1  g416(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n595_), .A2(new_n598_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n595_), .A2(KEYINPUT44), .A3(new_n598_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n571_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(G43gat), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n589_), .A2(G43gat), .A3(new_n419_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n618_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n618_), .ZN(new_n628_));
  AOI211_X1 g427(.A(new_n625_), .B(new_n628_), .C1(new_n623_), .C2(G43gat), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1330gat));
  NAND2_X1  g429(.A1(new_n601_), .A2(new_n579_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G50gat), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n470_), .A2(G50gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT106), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n632_), .B1(new_n589_), .B2(new_n634_), .ZN(G1331gat));
  INV_X1    g434(.A(G57gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n542_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n523_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n306_), .A2(new_n327_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n278_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n640_), .B2(new_n507_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT107), .Z(new_n642_));
  INV_X1    g441(.A(new_n543_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n278_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n327_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n551_), .A2(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n646_), .A2(new_n636_), .A3(new_n507_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n642_), .A2(new_n647_), .ZN(G1332gat));
  OAI21_X1  g447(.A(G64gat), .B1(new_n646_), .B2(new_n505_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT48), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n505_), .A2(G64gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n640_), .B2(new_n651_), .ZN(G1333gat));
  OAI21_X1  g451(.A(G71gat), .B1(new_n646_), .B2(new_n419_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n419_), .A2(G71gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n640_), .B2(new_n656_), .ZN(G1334gat));
  OR3_X1    g456(.A1(new_n640_), .A2(G78gat), .A3(new_n470_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n551_), .A2(new_n579_), .A3(new_n645_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT50), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n660_), .A3(G78gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n659_), .B2(G78gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT109), .ZN(G1335gat));
  NOR2_X1   g464(.A1(new_n644_), .A2(new_n587_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n638_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n219_), .A3(new_n383_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n278_), .A2(new_n542_), .A3(new_n327_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n383_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n669_), .B1(new_n672_), .B2(new_n219_), .ZN(G1336gat));
  NAND3_X1  g472(.A1(new_n668_), .A2(new_n220_), .A3(new_n504_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n671_), .A2(new_n504_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(new_n220_), .ZN(G1337gat));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n571_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n668_), .A2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n671_), .A2(new_n571_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n677_), .B(new_n679_), .C1(new_n680_), .C2(new_n234_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g481(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI211_X1 g483(.A(KEYINPUT111), .B(new_n216_), .C1(new_n671_), .C2(new_n579_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT111), .ZN(new_n686_));
  INV_X1    g485(.A(new_n670_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n506_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n470_), .A2(new_n504_), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n689_), .A2(new_n507_), .B1(new_n520_), .B2(new_n470_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n690_), .B2(new_n571_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n592_), .B1(new_n691_), .B2(new_n306_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n594_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n579_), .B(new_n687_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n686_), .B1(new_n694_), .B2(G106gat), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT52), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n685_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n470_), .A2(G106gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n668_), .A2(new_n698_), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n470_), .B(new_n670_), .C1(new_n591_), .C2(new_n594_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT111), .B1(new_n700_), .B2(new_n216_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n701_), .B2(KEYINPUT52), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n684_), .B1(new_n697_), .B2(new_n702_), .ZN(new_n703_));
  AOI22_X1  g502(.A1(new_n695_), .A2(new_n696_), .B1(new_n668_), .B2(new_n698_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(KEYINPUT52), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n704_), .B(new_n683_), .C1(new_n705_), .C2(new_n685_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1339gat));
  INV_X1    g506(.A(KEYINPUT120), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT113), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n328_), .A2(new_n543_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(KEYINPUT54), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT54), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n328_), .A2(KEYINPUT113), .A3(new_n712_), .A4(new_n543_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(KEYINPUT54), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n711_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n550_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n716_), .A2(KEYINPUT57), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n524_), .A2(new_n525_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n528_), .A2(new_n529_), .A3(new_n526_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n535_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n537_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n275_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n274_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n270_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n637_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n242_), .A2(new_n251_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT114), .B1(new_n268_), .B2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n259_), .B1(new_n249_), .B2(new_n209_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n730_), .B1(new_n287_), .B2(new_n266_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT114), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n252_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n258_), .B1(new_n729_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT115), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n731_), .B2(new_n252_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n265_), .A2(new_n267_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n728_), .A2(new_n738_), .A3(KEYINPUT114), .A4(new_n730_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(KEYINPUT115), .A3(new_n258_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(new_n730_), .A3(new_n269_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT116), .B1(new_n742_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n748_), .B(new_n745_), .C1(new_n736_), .C2(new_n741_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n274_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT115), .B1(new_n740_), .B2(new_n258_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n735_), .B(new_n257_), .C1(new_n737_), .C2(new_n739_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n746_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n748_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n746_), .B(KEYINPUT116), .C1(new_n753_), .C2(new_n754_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(KEYINPUT56), .A3(new_n274_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n727_), .B1(new_n752_), .B2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n724_), .B1(new_n760_), .B2(KEYINPUT117), .ZN(new_n761_));
  INV_X1    g560(.A(new_n727_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT56), .B1(new_n758_), .B2(new_n274_), .ZN(new_n763_));
  AOI211_X1 g562(.A(new_n751_), .B(new_n725_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n717_), .B1(new_n761_), .B2(new_n767_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n726_), .B(new_n721_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n305_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n726_), .A2(new_n721_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n752_), .B2(new_n759_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n771_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n723_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n760_), .A2(KEYINPUT117), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n550_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n768_), .B(new_n775_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n715_), .B1(new_n780_), .B2(new_n327_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n579_), .A2(new_n504_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n507_), .A2(new_n419_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n784_), .A2(KEYINPUT59), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n708_), .B1(new_n781_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n776_), .A2(new_n777_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n788_), .A2(new_n717_), .B1(new_n774_), .B2(new_n771_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n716_), .B1(new_n761_), .B2(new_n767_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n779_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n553_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT120), .B(new_n785_), .C1(new_n793_), .C2(new_n715_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n306_), .B1(new_n773_), .B2(KEYINPUT58), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n769_), .A2(new_n770_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT119), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n771_), .A2(new_n799_), .A3(new_n774_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(new_n792_), .A3(new_n768_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n715_), .B1(new_n802_), .B2(new_n327_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT59), .B1(new_n803_), .B2(new_n784_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n795_), .A2(new_n643_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(G113gat), .ZN(new_n806_));
  INV_X1    g605(.A(new_n784_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n790_), .A2(new_n791_), .B1(new_n788_), .B2(new_n717_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n553_), .B1(new_n808_), .B2(new_n801_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n807_), .B1(new_n809_), .B2(new_n715_), .ZN(new_n810_));
  OR3_X1    g609(.A1(new_n810_), .A2(G113gat), .A3(new_n542_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n806_), .A2(new_n811_), .ZN(G1340gat));
  NAND3_X1  g611(.A1(new_n795_), .A2(new_n278_), .A3(new_n804_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G120gat), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT60), .ZN(new_n815_));
  AOI21_X1  g614(.A(G120gat), .B1(new_n278_), .B2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT121), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n815_), .B2(G120gat), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n807_), .B(new_n818_), .C1(new_n809_), .C2(new_n715_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT122), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n814_), .A2(new_n821_), .ZN(G1341gat));
  NAND3_X1  g621(.A1(new_n795_), .A2(new_n553_), .A3(new_n804_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G127gat), .ZN(new_n824_));
  OR3_X1    g623(.A1(new_n810_), .A2(G127gat), .A3(new_n327_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1342gat));
  INV_X1    g625(.A(G134gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n810_), .B2(new_n716_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT123), .B(new_n827_), .C1(new_n810_), .C2(new_n716_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n787_), .A2(new_n794_), .B1(new_n810_), .B2(KEYINPUT59), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n305_), .A2(new_n827_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n830_), .A2(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(G1343gat));
  NOR2_X1   g633(.A1(new_n803_), .A2(new_n571_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n470_), .A2(new_n507_), .A3(new_n504_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G141gat), .B1(new_n837_), .B2(new_n542_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n835_), .A2(new_n343_), .A3(new_n637_), .A4(new_n836_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1344gat));
  OAI21_X1  g639(.A(G148gat), .B1(new_n837_), .B2(new_n644_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n835_), .A2(new_n344_), .A3(new_n278_), .A4(new_n836_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1345gat));
  XNOR2_X1  g642(.A(KEYINPUT61), .B(G155gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n837_), .B2(new_n327_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n844_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n835_), .A2(new_n553_), .A3(new_n836_), .A4(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1346gat));
  OAI21_X1  g647(.A(G162gat), .B1(new_n837_), .B2(new_n305_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n835_), .A2(new_n353_), .A3(new_n550_), .A4(new_n836_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1347gat));
  NAND2_X1  g650(.A1(new_n420_), .A2(new_n504_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT124), .Z(new_n853_));
  OR3_X1    g652(.A1(new_n853_), .A2(new_n579_), .A3(new_n542_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n781_), .A2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n477_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n855_), .B2(G169gat), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n855_), .A2(new_n857_), .A3(G169gat), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n781_), .A2(new_n854_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT125), .B1(new_n862_), .B2(new_n387_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n863_), .A3(KEYINPUT62), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n864_), .ZN(G1348gat));
  NOR3_X1   g664(.A1(new_n781_), .A2(new_n579_), .A3(new_n853_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G176gat), .B1(new_n866_), .B2(new_n278_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n803_), .A2(new_n579_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n853_), .A2(new_n388_), .A3(new_n644_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(G1349gat));
  NOR2_X1   g669(.A1(new_n853_), .A2(new_n327_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G183gat), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n327_), .A2(new_n472_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n866_), .B2(new_n873_), .ZN(G1350gat));
  NAND2_X1  g673(.A1(new_n866_), .A2(new_n306_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G190gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n866_), .A2(new_n392_), .A3(new_n550_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1351gat));
  NOR3_X1   g677(.A1(new_n470_), .A2(new_n383_), .A3(new_n505_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n419_), .B(new_n879_), .C1(new_n809_), .C2(new_n715_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(G197gat), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n880_), .A2(new_n542_), .A3(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n835_), .A2(new_n637_), .A3(new_n879_), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT126), .B(G197gat), .Z(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1352gat));
  NOR2_X1   g685(.A1(new_n880_), .A2(new_n644_), .ZN(new_n887_));
  INV_X1    g686(.A(G204gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1353gat));
  AOI21_X1  g688(.A(new_n327_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n890_));
  XOR2_X1   g689(.A(new_n890_), .B(KEYINPUT127), .Z(new_n891_));
  NOR2_X1   g690(.A1(new_n880_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1354gat));
  OAI21_X1  g693(.A(G218gat), .B1(new_n880_), .B2(new_n305_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n716_), .A2(G218gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n880_), .B2(new_n896_), .ZN(G1355gat));
endmodule


