//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT77), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G169gat), .B(G197gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G229gat), .A2(G233gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G29gat), .B(G36gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217_));
  INV_X1    g016(.A(G1gat), .ZN(new_n218_));
  INV_X1    g017(.A(G8gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT14), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G1gat), .B(G8gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT75), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n211_), .A2(KEYINPUT15), .A3(new_n213_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n216_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n221_), .B(new_n222_), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n214_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n216_), .A2(new_n225_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT75), .B1(new_n230_), .B2(new_n227_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n207_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n223_), .B(new_n214_), .Z(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(new_n206_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n205_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT78), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n237_), .B(new_n205_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  OR3_X1    g038(.A1(new_n232_), .A2(new_n234_), .A3(KEYINPUT76), .ZN(new_n240_));
  INV_X1    g039(.A(new_n205_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT76), .B1(new_n232_), .B2(new_n234_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(G141gat), .A2(G148gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G155gat), .A2(G162gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT1), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT83), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n252_), .A2(G155gat), .A3(G162gat), .ZN(new_n253_));
  INV_X1    g052(.A(G155gat), .ZN(new_n254_));
  INV_X1    g053(.A(G162gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT83), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n251_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT84), .B1(new_n250_), .B2(KEYINPUT1), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT84), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(G155gat), .A4(G162gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n249_), .B1(new_n257_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT29), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n248_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n246_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n254_), .A2(new_n255_), .A3(KEYINPUT83), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n252_), .B1(G155gat), .B2(G162gat), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n272_), .A2(new_n273_), .B1(G155gat), .B2(G162gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n263_), .A2(new_n264_), .A3(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(KEYINPUT28), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT28), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G22gat), .B(G50gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G78gat), .B(G106gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G228gat), .A2(G233gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT87), .ZN(new_n284_));
  INV_X1    g083(.A(G197gat), .ZN(new_n285_));
  INV_X1    g084(.A(G204gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G197gat), .A2(G204gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT21), .A3(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(G197gat), .A2(G204gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G197gat), .A2(G204gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n289_), .B(new_n290_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT86), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT21), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n299_), .A2(KEYINPUT85), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(KEYINPUT85), .ZN(new_n301_));
  OAI22_X1  g100(.A1(new_n300_), .A2(new_n301_), .B1(new_n292_), .B2(new_n291_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n302_), .A2(new_n296_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n284_), .B1(new_n298_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n249_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n258_), .A2(new_n261_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n272_), .A2(new_n273_), .B1(KEYINPUT1), .B2(new_n250_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n271_), .A2(new_n274_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT29), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n283_), .A2(KEYINPUT87), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n304_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n304_), .B2(new_n310_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n282_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n277_), .A2(new_n278_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n279_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n298_), .A2(new_n303_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n264_), .B1(new_n263_), .B2(new_n275_), .ZN(new_n319_));
  OAI211_X1 g118(.A(KEYINPUT87), .B(new_n283_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n304_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n281_), .ZN(new_n322_));
  AND4_X1   g121(.A1(new_n280_), .A2(new_n314_), .A3(new_n317_), .A4(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n314_), .A2(KEYINPUT88), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n320_), .A2(new_n321_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT88), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n282_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n325_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n317_), .A2(new_n280_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n330_), .A2(KEYINPUT89), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT89), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n328_), .B1(new_n327_), .B2(new_n282_), .ZN(new_n335_));
  AOI211_X1 g134(.A(KEYINPUT88), .B(new_n281_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n322_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n337_), .B2(new_n331_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n324_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT90), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT89), .B1(new_n330_), .B2(new_n332_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n334_), .A3(new_n331_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT90), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n324_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G8gat), .B(G36gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT18), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT25), .B1(KEYINPUT79), .B2(G183gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n355_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n360_), .A3(G183gat), .ZN(new_n361_));
  INV_X1    g160(.A(G190gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT26), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT26), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G190gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT81), .B1(new_n359_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(G169gat), .ZN(new_n368_));
  INV_X1    g167(.A(G176gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(KEYINPUT24), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT23), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(G183gat), .A3(G190gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  OR3_X1    g176(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n372_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n380_));
  INV_X1    g179(.A(G183gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n382_), .B(KEYINPUT25), .C1(KEYINPUT80), .C2(new_n356_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n363_), .A2(new_n365_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .A4(new_n361_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n367_), .A2(new_n379_), .A3(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G169gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n382_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n390_), .A2(G190gat), .A3(new_n357_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n373_), .B(new_n375_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n389_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n387_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n354_), .B1(new_n394_), .B2(new_n318_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT22), .B(G169gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n369_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n371_), .B(KEYINPUT91), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT92), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT92), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G183gat), .A2(G190gat), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n392_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT25), .B(G183gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n384_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n379_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n298_), .A2(new_n303_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n353_), .B1(new_n395_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n318_), .A2(new_n408_), .A3(new_n405_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n387_), .A2(new_n393_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n410_), .ZN(new_n415_));
  AND4_X1   g214(.A1(KEYINPUT20), .A2(new_n413_), .A3(new_n415_), .A4(new_n353_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n350_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n415_), .A3(KEYINPUT20), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n352_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n395_), .A2(new_n353_), .A3(new_n411_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT32), .A4(new_n349_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT94), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G127gat), .B(G134gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G113gat), .B(G120gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n426_), .A2(new_n427_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT95), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n430_), .B(new_n431_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n263_), .B(new_n275_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT4), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n263_), .A2(new_n275_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n435_), .A2(new_n431_), .A3(new_n436_), .A4(new_n430_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n425_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT97), .ZN(new_n441_));
  XOR2_X1   g240(.A(G1gat), .B(G29gat), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n441_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G57gat), .B(G85gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n435_), .A2(new_n430_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n424_), .B1(new_n447_), .B2(new_n433_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n439_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n445_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n444_), .B(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n438_), .B2(new_n448_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(new_n453_), .A3(KEYINPUT99), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT99), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n439_), .A2(new_n446_), .A3(new_n455_), .A4(new_n449_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n422_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n457_), .A2(KEYINPUT100), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n434_), .A2(new_n425_), .A3(new_n437_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n447_), .A2(new_n424_), .A3(new_n433_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n446_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n461_), .B1(new_n453_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n349_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n318_), .B1(new_n408_), .B2(new_n405_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n410_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n352_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n468_), .B(new_n349_), .C1(new_n352_), .C2(new_n418_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT93), .B(new_n464_), .C1(new_n412_), .C2(new_n416_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n463_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n453_), .A2(new_n462_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT98), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT98), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n453_), .A2(new_n476_), .A3(new_n462_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n473_), .A2(new_n478_), .B1(new_n457_), .B2(KEYINPUT100), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n340_), .A2(new_n345_), .A3(new_n458_), .A4(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT27), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n471_), .A2(new_n481_), .A3(new_n472_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n419_), .A2(new_n420_), .ZN(new_n483_));
  OAI211_X1 g282(.A(KEYINPUT27), .B(new_n469_), .C1(new_n483_), .C2(new_n349_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n454_), .A2(new_n456_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n344_), .B1(new_n343_), .B2(new_n324_), .ZN(new_n487_));
  AOI211_X1 g286(.A(KEYINPUT90), .B(new_n323_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G71gat), .B(G99gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT82), .B(G43gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n414_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(new_n430_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G227gat), .A2(G233gat), .ZN(new_n495_));
  INV_X1    g294(.A(G15gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT30), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT31), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n494_), .B(new_n499_), .Z(new_n500_));
  NAND3_X1  g299(.A1(new_n480_), .A2(new_n489_), .A3(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n487_), .A2(new_n488_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n482_), .A2(new_n484_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n485_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n245_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT12), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT6), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT9), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(G85gat), .A3(G92gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G85gat), .B(G92gat), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n510_), .B(new_n512_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT64), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n517_), .B2(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(G106gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(KEYINPUT64), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n514_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n523_));
  INV_X1    g322(.A(G99gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n519_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT65), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n523_), .A2(new_n524_), .A3(new_n519_), .A4(KEYINPUT65), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n510_), .A2(new_n522_), .A3(new_n527_), .A4(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n513_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT8), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT8), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n533_), .A3(new_n530_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n521_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT66), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(KEYINPUT66), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G71gat), .B(G78gat), .ZN(new_n542_));
  OAI22_X1  g341(.A1(new_n538_), .A2(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n538_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n541_), .A2(new_n542_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n539_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n508_), .B1(new_n535_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n535_), .A2(new_n547_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n521_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n534_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT67), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n533_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT67), .B1(new_n532_), .B2(new_n534_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n551_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n547_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(KEYINPUT12), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n550_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n549_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n535_), .A2(new_n547_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G120gat), .B(G148gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G176gat), .B(G204gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n561_), .A2(new_n565_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n575_), .B1(new_n578_), .B2(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT37), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n535_), .B2(new_n214_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n585_), .B1(new_n587_), .B2(KEYINPUT71), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n553_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n532_), .A2(KEYINPUT67), .A3(new_n534_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n521_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n587_), .B1(new_n591_), .B2(new_n230_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n592_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT72), .ZN(new_n597_));
  XOR2_X1   g396(.A(G134gat), .B(G162gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT36), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n581_), .B1(new_n595_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n593_), .A2(KEYINPUT73), .A3(new_n594_), .A4(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n593_), .A2(new_n594_), .A3(new_n604_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT73), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT74), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n595_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n593_), .A2(KEYINPUT74), .A3(new_n594_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n600_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n607_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n610_), .B1(new_n616_), .B2(KEYINPUT37), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n223_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n547_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT16), .ZN(new_n623_));
  XOR2_X1   g422(.A(G183gat), .B(G211gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n620_), .A2(new_n621_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(KEYINPUT17), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n620_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n617_), .A2(new_n630_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n507_), .A2(new_n580_), .A3(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n218_), .A3(new_n504_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n616_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n636_));
  AND4_X1   g435(.A1(new_n244_), .A2(new_n636_), .A3(new_n580_), .A4(new_n629_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n218_), .B1(new_n637_), .B2(new_n504_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n634_), .B2(new_n633_), .ZN(G1324gat));
  INV_X1    g439(.A(new_n503_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n219_), .B1(new_n637_), .B2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT39), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n632_), .A2(new_n219_), .A3(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g445(.A(new_n500_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n496_), .B1(new_n637_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT41), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n632_), .A2(new_n496_), .A3(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n502_), .B(KEYINPUT101), .Z(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n637_), .B2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT42), .Z(new_n656_));
  NAND3_X1  g455(.A1(new_n632_), .A2(new_n654_), .A3(new_n652_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1327gat));
  NAND2_X1  g457(.A1(new_n616_), .A2(new_n630_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT104), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n507_), .A3(new_n580_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n660_), .A2(KEYINPUT105), .A3(new_n507_), .A4(new_n580_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n665_), .A2(G29gat), .A3(new_n485_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n501_), .A2(new_n506_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n617_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n667_), .A2(KEYINPUT102), .A3(new_n668_), .A4(new_n617_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n667_), .A2(new_n617_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT43), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n580_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n676_), .A2(new_n245_), .A3(new_n629_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n504_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n680_), .A2(new_n681_), .A3(G29gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n680_), .B2(G29gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n666_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  INV_X1    g483(.A(G36gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n679_), .B2(new_n641_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n503_), .B(KEYINPUT106), .Z(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(G36gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n663_), .A2(new_n664_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT107), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n663_), .A2(new_n692_), .A3(new_n664_), .A4(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT45), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n687_), .A2(KEYINPUT46), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n694_), .B(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n699_), .B2(new_n686_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n696_), .A2(new_n700_), .ZN(G1329gat));
  NAND3_X1  g500(.A1(new_n679_), .A2(G43gat), .A3(new_n647_), .ZN(new_n702_));
  INV_X1    g501(.A(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n665_), .B2(new_n500_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(G1330gat));
  INV_X1    g506(.A(G50gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n502_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n663_), .A2(new_n654_), .A3(new_n664_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n679_), .A2(new_n709_), .B1(new_n708_), .B2(new_n710_), .ZN(G1331gat));
  NOR3_X1   g510(.A1(new_n580_), .A2(new_n244_), .A3(new_n630_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n636_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n485_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n244_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n716_), .A2(new_n676_), .A3(new_n631_), .ZN(new_n717_));
  INV_X1    g516(.A(G57gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n504_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n719_), .ZN(G1332gat));
  INV_X1    g519(.A(G64gat), .ZN(new_n721_));
  INV_X1    g520(.A(new_n688_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n713_), .B2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT48), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n717_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT109), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n713_), .B2(new_n647_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT49), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n717_), .A2(new_n728_), .A3(new_n647_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT110), .Z(G1334gat));
  INV_X1    g532(.A(G78gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n713_), .B2(new_n654_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT50), .Z(new_n736_));
  NAND3_X1  g535(.A1(new_n717_), .A2(new_n654_), .A3(new_n734_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1335gat));
  NOR3_X1   g537(.A1(new_n580_), .A2(new_n244_), .A3(new_n629_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n675_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n485_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n660_), .A2(new_n676_), .A3(new_n716_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT111), .ZN(new_n744_));
  INV_X1    g543(.A(G85gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n504_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n742_), .A2(new_n746_), .ZN(G1336gat));
  OAI21_X1  g546(.A(G92gat), .B1(new_n741_), .B2(new_n688_), .ZN(new_n748_));
  INV_X1    g547(.A(G92gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n744_), .A2(new_n749_), .A3(new_n641_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1337gat));
  AOI21_X1  g550(.A(new_n524_), .B1(new_n740_), .B2(new_n647_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n500_), .A2(new_n517_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n744_), .B2(new_n753_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g554(.A(new_n502_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n744_), .A2(new_n519_), .A3(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n675_), .A2(new_n756_), .A3(new_n739_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(G106gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT113), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n758_), .A2(new_n763_), .A3(new_n760_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n759_), .B1(new_n758_), .B2(G106gat), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n762_), .B(new_n764_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n766_), .A2(new_n765_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n757_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT53), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n757_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT122), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n244_), .A2(new_n574_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n560_), .B1(new_n550_), .B2(new_n559_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n561_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n558_), .A2(KEYINPUT12), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n549_), .B(new_n548_), .C1(new_n591_), .C2(new_n780_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n781_), .A2(new_n778_), .A3(new_n562_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n779_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(KEYINPUT56), .A4(new_n571_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n778_), .B1(new_n781_), .B2(new_n562_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n781_), .A2(new_n562_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(KEYINPUT56), .B(new_n571_), .C1(new_n789_), .C2(new_n782_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT116), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT56), .B1(new_n784_), .B2(new_n571_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n776_), .B(new_n786_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n229_), .A2(new_n231_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n206_), .B1(new_n794_), .B2(KEYINPUT117), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(KEYINPUT117), .B2(new_n794_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n205_), .B1(new_n233_), .B2(new_n206_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n236_), .A2(new_n238_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(new_n574_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n573_), .B1(new_n561_), .B2(new_n565_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n798_), .B(new_n799_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n799_), .B1(new_n575_), .B2(new_n798_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n616_), .B1(new_n793_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT119), .B1(new_n806_), .B2(KEYINPUT57), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n798_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT118), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n802_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n776_), .A2(new_n786_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n571_), .B1(new_n789_), .B2(new_n782_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(KEYINPUT116), .A3(new_n790_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n812_), .B1(new_n813_), .B2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n808_), .B(new_n809_), .C1(new_n818_), .C2(new_n616_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n807_), .A2(new_n819_), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n615_), .A2(new_n581_), .B1(new_n606_), .B2(new_n609_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n790_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n784_), .A2(KEYINPUT120), .A3(KEYINPUT56), .A4(new_n571_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n816_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n798_), .A2(new_n574_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT121), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n821_), .B1(new_n828_), .B2(KEYINPUT58), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n829_), .A2(new_n833_), .B1(KEYINPUT57), .B2(new_n806_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n629_), .B1(new_n820_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n631_), .A2(new_n245_), .A3(new_n580_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n631_), .A2(new_n245_), .A3(new_n580_), .A4(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n774_), .B1(new_n835_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n806_), .A2(KEYINPUT57), .ZN(new_n844_));
  INV_X1    g643(.A(new_n833_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n617_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n807_), .A2(new_n819_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n630_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT122), .A3(new_n841_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n843_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n756_), .A2(new_n641_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n504_), .A3(new_n647_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(G113gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n244_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n853_), .A2(KEYINPUT59), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n806_), .A2(KEYINPUT57), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n630_), .B1(new_n847_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n842_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n859_), .A2(new_n860_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n857_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n849_), .A2(KEYINPUT122), .A3(new_n841_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT122), .B1(new_n849_), .B2(new_n841_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n853_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI211_X1 g667(.A(new_n245_), .B(new_n863_), .C1(new_n868_), .C2(KEYINPUT59), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n856_), .B1(new_n869_), .B2(new_n855_), .ZN(G1340gat));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n580_), .A2(KEYINPUT60), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT124), .B(G120gat), .ZN(new_n873_));
  MUX2_X1   g672(.A(KEYINPUT60), .B(new_n872_), .S(new_n873_), .Z(new_n874_));
  NAND3_X1  g673(.A1(new_n854_), .A2(new_n871_), .A3(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n866_), .A2(new_n867_), .A3(new_n874_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT125), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n580_), .B(new_n863_), .C1(new_n868_), .C2(KEYINPUT59), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n873_), .ZN(G1341gat));
  INV_X1    g679(.A(G127gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n854_), .A2(new_n881_), .A3(new_n629_), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n630_), .B(new_n863_), .C1(new_n868_), .C2(KEYINPUT59), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1342gat));
  INV_X1    g683(.A(G134gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n854_), .A2(new_n885_), .A3(new_n616_), .ZN(new_n886_));
  AOI211_X1 g685(.A(new_n821_), .B(new_n863_), .C1(new_n868_), .C2(KEYINPUT59), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1343gat));
  NOR3_X1   g687(.A1(new_n722_), .A2(new_n485_), .A3(new_n647_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n843_), .A2(new_n756_), .A3(new_n850_), .A4(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n245_), .ZN(new_n891_));
  XOR2_X1   g690(.A(new_n891_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n580_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g693(.A1(new_n890_), .A2(new_n630_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n895_), .B(new_n896_), .Z(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n890_), .B2(new_n821_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n615_), .A2(G162gat), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n866_), .A2(new_n756_), .A3(new_n889_), .A4(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(KEYINPUT126), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n898_), .A2(new_n903_), .A3(new_n900_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1347gat));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n861_), .A2(new_n862_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n722_), .A2(new_n505_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n654_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n245_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n906_), .B1(new_n911_), .B2(new_n368_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n396_), .ZN(new_n913_));
  OAI211_X1 g712(.A(KEYINPUT62), .B(G169gat), .C1(new_n910_), .C2(new_n245_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(G1348gat));
  INV_X1    g714(.A(new_n910_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G176gat), .B1(new_n916_), .B2(new_n676_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n851_), .A2(new_n756_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n908_), .A2(new_n369_), .A3(new_n580_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n918_), .B2(new_n919_), .ZN(G1349gat));
  NOR3_X1   g719(.A1(new_n910_), .A2(new_n406_), .A3(new_n630_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n918_), .A2(new_n505_), .A3(new_n629_), .A4(new_n722_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n390_), .A2(new_n357_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n910_), .B2(new_n821_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n616_), .A2(new_n384_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n910_), .B2(new_n926_), .ZN(G1351gat));
  NOR3_X1   g726(.A1(new_n688_), .A2(new_n504_), .A3(new_n647_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n843_), .A2(new_n756_), .A3(new_n850_), .A4(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n245_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(new_n285_), .ZN(G1352gat));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n580_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n286_), .ZN(G1353gat));
  NOR2_X1   g732(.A1(new_n929_), .A2(new_n630_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n934_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT63), .B(G211gat), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n929_), .A2(new_n630_), .A3(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n935_), .A2(new_n937_), .ZN(G1354gat));
  INV_X1    g737(.A(G218gat), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n929_), .A2(new_n939_), .A3(new_n821_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n929_), .A2(new_n615_), .ZN(new_n941_));
  AOI21_X1  g740(.A(G218gat), .B1(new_n941_), .B2(KEYINPUT127), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n929_), .B2(new_n615_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n940_), .B1(new_n942_), .B2(new_n944_), .ZN(G1355gat));
endmodule


