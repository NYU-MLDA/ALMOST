//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(KEYINPUT82), .A3(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT21), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n210_), .B2(new_n205_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n211_), .A2(KEYINPUT83), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(KEYINPUT83), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n206_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n205_), .A2(new_n202_), .A3(new_n204_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(G141gat), .ZN(new_n219_));
  INV_X1    g018(.A(G148gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT1), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n218_), .B(new_n221_), .C1(new_n224_), .C2(new_n226_), .ZN(new_n227_));
  OR3_X1    g026(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n222_), .B(KEYINPUT78), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n225_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n217_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT81), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n236_), .A2(KEYINPUT80), .A3(KEYINPUT29), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n241_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT84), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n242_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT85), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n251_), .A2(KEYINPUT86), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT86), .B1(new_n251_), .B2(new_n254_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n253_), .B(new_n242_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT79), .B(KEYINPUT28), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G22gat), .B(G50gat), .Z(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(new_n236_), .B2(KEYINPUT29), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n267_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n255_), .A2(new_n256_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n251_), .A2(new_n252_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n267_), .B1(new_n270_), .B2(new_n257_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT87), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G226gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT19), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT23), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(G183gat), .B2(G190gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(G183gat), .A3(G190gat), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G169gat), .ZN(new_n286_));
  INV_X1    g085(.A(G176gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(KEYINPUT26), .B(G190gat), .Z(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT25), .B(G183gat), .Z(new_n290_));
  OAI211_X1 g089(.A(new_n283_), .B(new_n288_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(G169gat), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n280_), .A2(KEYINPUT75), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n280_), .A2(KEYINPUT75), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n278_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n293_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n276_), .B1(new_n217_), .B2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n211_), .B(KEYINPUT83), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n215_), .B1(new_n301_), .B2(new_n206_), .ZN(new_n302_));
  OR3_X1    g101(.A1(new_n296_), .A2(KEYINPUT76), .A3(new_n282_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT76), .B1(new_n296_), .B2(new_n282_), .ZN(new_n304_));
  INV_X1    g103(.A(G190gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT74), .B1(new_n305_), .B2(KEYINPUT26), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n290_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n289_), .A2(KEYINPUT74), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n309_), .A2(new_n288_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n303_), .A2(new_n304_), .A3(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n293_), .B1(new_n281_), .B2(new_n297_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n302_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n275_), .B1(new_n300_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n291_), .A2(new_n298_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n276_), .B1(new_n316_), .B2(new_n302_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n312_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n217_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n319_), .A3(new_n275_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G8gat), .B(G36gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n315_), .A2(new_n320_), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n275_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n300_), .A2(new_n275_), .A3(new_n313_), .ZN(new_n330_));
  OAI211_X1 g129(.A(KEYINPUT32), .B(new_n326_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT77), .ZN(new_n339_));
  XOR2_X1   g138(.A(G113gat), .B(G120gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(new_n236_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n236_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(KEYINPUT4), .A3(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT89), .B(KEYINPUT4), .Z(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n236_), .A3(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n346_), .A2(KEYINPUT90), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(KEYINPUT90), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n344_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n337_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  AOI211_X1 g154(.A(new_n336_), .B(new_n353_), .C1(new_n349_), .C2(new_n351_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n328_), .B(new_n331_), .C1(new_n355_), .C2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n346_), .B(KEYINPUT90), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n350_), .B1(new_n358_), .B2(new_n344_), .ZN(new_n359_));
  OAI211_X1 g158(.A(KEYINPUT33), .B(new_n336_), .C1(new_n359_), .C2(new_n353_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n350_), .A3(new_n344_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n342_), .A2(new_n343_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n336_), .B1(new_n363_), .B2(new_n351_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n361_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n360_), .B1(new_n355_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n320_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n325_), .B1(new_n367_), .B2(new_n314_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n315_), .A2(new_n326_), .A3(new_n320_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n357_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n251_), .A2(new_n254_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n251_), .A2(KEYINPUT86), .A3(new_n254_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n374_), .A2(new_n257_), .A3(new_n267_), .A4(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT87), .ZN(new_n377_));
  INV_X1    g176(.A(new_n271_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n272_), .A2(new_n371_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT92), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT92), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n272_), .A2(new_n371_), .A3(new_n382_), .A4(new_n379_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n272_), .A2(new_n379_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n355_), .A2(new_n356_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT27), .B1(new_n368_), .B2(new_n369_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n325_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(new_n369_), .A3(KEYINPUT27), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n386_), .A2(new_n387_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n381_), .A2(new_n383_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT30), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n318_), .B(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n398_), .A2(new_n341_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n341_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G71gat), .B(G99gat), .ZN(new_n402_));
  INV_X1    g201(.A(G43gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT31), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n399_), .A2(new_n405_), .A3(new_n400_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT27), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n370_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(KEYINPUT93), .A3(new_n389_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT93), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n390_), .B2(new_n387_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n409_), .A2(new_n386_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n415_), .A2(new_n272_), .A3(new_n416_), .A4(new_n379_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT94), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n272_), .A2(new_n379_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n420_), .A2(KEYINPUT94), .A3(new_n415_), .A4(new_n416_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n393_), .A2(new_n409_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G113gat), .B(G141gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G169gat), .B(G197gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  NAND2_X1  g224(.A1(G229gat), .A2(G233gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G15gat), .B(G22gat), .ZN(new_n427_));
  INV_X1    g226(.A(G1gat), .ZN(new_n428_));
  INV_X1    g227(.A(G8gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT14), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G1gat), .B(G8gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G29gat), .B(G36gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G43gat), .B(G50gat), .Z(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G43gat), .B(G50gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n433_), .A2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n431_), .A2(new_n432_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n431_), .A2(new_n432_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n426_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n446_), .A2(KEYINPUT69), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(KEYINPUT69), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT15), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n440_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n437_), .A2(KEYINPUT15), .A3(new_n439_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n433_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT70), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n426_), .B(KEYINPUT71), .Z(new_n456_));
  AND2_X1   g255(.A1(new_n445_), .A2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  OAI211_X1 g257(.A(KEYINPUT72), .B(new_n425_), .C1(new_n449_), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n425_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n447_), .A2(new_n448_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT72), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n460_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT73), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n422_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G120gat), .B(G148gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT5), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G176gat), .B(G204gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G230gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  OR2_X1    g272(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G85gat), .ZN(new_n478_));
  INV_X1    g277(.A(G92gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G85gat), .A2(G92gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(KEYINPUT9), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT9), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n486_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n473_), .B1(new_n483_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n493_), .A2(new_n494_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n495_), .A2(KEYINPUT64), .A3(new_n482_), .A4(new_n477_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498_));
  INV_X1    g297(.A(G99gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n475_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT7), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n493_), .A2(new_n494_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT7), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n498_), .A2(new_n503_), .A3(new_n499_), .A4(new_n475_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n501_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n480_), .A2(new_n481_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT8), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(KEYINPUT8), .A3(new_n506_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G71gat), .B(G78gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(KEYINPUT11), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n514_));
  INV_X1    g313(.A(new_n512_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n513_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n497_), .A2(new_n509_), .A3(new_n510_), .A4(new_n518_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n492_), .A2(new_n496_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n520_), .B2(new_n510_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n521_), .B2(KEYINPUT66), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n497_), .A2(new_n510_), .A3(new_n509_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n518_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n523_), .A2(KEYINPUT66), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n472_), .B1(new_n522_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n472_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n524_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(KEYINPUT12), .A3(new_n519_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n523_), .A2(new_n531_), .A3(new_n524_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n528_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n527_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n519_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(new_n529_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n528_), .B1(new_n538_), .B2(new_n525_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT67), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n471_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n519_), .A2(KEYINPUT12), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(new_n521_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n532_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n472_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n539_), .A2(KEYINPUT67), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n527_), .A2(new_n534_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n470_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n541_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n549_), .A2(KEYINPUT13), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(KEYINPUT13), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n451_), .A2(new_n452_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n523_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n520_), .A2(new_n441_), .A3(new_n510_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT68), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n557_), .A2(new_n561_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G134gat), .B(G162gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n570_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n567_), .A2(new_n569_), .A3(new_n574_), .A4(new_n573_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n577_), .A2(KEYINPUT37), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT37), .B1(new_n577_), .B2(new_n578_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n433_), .B(new_n518_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  OR3_X1    g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(KEYINPUT17), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n582_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n466_), .A2(new_n552_), .A3(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n597_), .A2(G1gat), .A3(new_n385_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n598_), .A2(KEYINPUT38), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(KEYINPUT38), .ZN(new_n600_));
  INV_X1    g399(.A(new_n552_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(new_n464_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n595_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT95), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n577_), .A2(new_n578_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n422_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n610_), .B2(new_n385_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n599_), .A2(new_n600_), .A3(new_n611_), .ZN(G1324gat));
  OAI21_X1  g411(.A(G8gat), .B1(new_n610_), .B2(new_n415_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT39), .ZN(new_n614_));
  INV_X1    g413(.A(new_n597_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n415_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n429_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(G1325gat));
  OAI21_X1  g419(.A(G15gat), .B1(new_n610_), .B2(new_n409_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT41), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n409_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n615_), .A2(new_n395_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(G1326gat));
  OR3_X1    g427(.A1(new_n597_), .A2(G22gat), .A3(new_n420_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n605_), .A2(new_n384_), .A3(new_n609_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT98), .B(KEYINPUT42), .Z(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(G22gat), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n630_), .B2(G22gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n629_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT99), .Z(G1327gat));
  NAND2_X1  g435(.A1(new_n608_), .A2(new_n595_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n601_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n465_), .ZN(new_n641_));
  AOI22_X1  g440(.A1(new_n380_), .A2(KEYINPUT92), .B1(new_n384_), .B2(new_n391_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n624_), .B1(new_n642_), .B2(new_n383_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n419_), .A2(new_n421_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n640_), .B(new_n641_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(G29gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n386_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n649_), .B1(new_n422_), .B2(new_n581_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT43), .B(new_n582_), .C1(new_n644_), .C2(new_n643_), .ZN(new_n651_));
  AND4_X1   g450(.A1(new_n595_), .A2(new_n650_), .A3(new_n602_), .A4(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(KEYINPUT100), .A3(KEYINPUT44), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n650_), .A2(new_n651_), .A3(new_n595_), .A4(new_n602_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n653_), .A2(new_n657_), .B1(new_n656_), .B2(new_n655_), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT101), .B(new_n647_), .C1(new_n658_), .C2(new_n386_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n653_), .A2(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n655_), .A2(new_n656_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n386_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n660_), .B1(new_n663_), .B2(G29gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n648_), .B1(new_n659_), .B2(new_n664_), .ZN(G1328gat));
  XNOR2_X1  g464(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n415_), .A2(G36gat), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT103), .B1(new_n645_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n466_), .A2(new_n671_), .A3(new_n640_), .A4(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT45), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n670_), .A2(KEYINPUT45), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n415_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT100), .B1(new_n652_), .B2(KEYINPUT44), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n655_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n677_), .B1(new_n681_), .B2(G36gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n667_), .B1(new_n682_), .B2(KEYINPUT104), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684_));
  INV_X1    g483(.A(G36gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n661_), .B2(new_n678_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n684_), .B(new_n666_), .C1(new_n686_), .C2(new_n677_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n687_), .ZN(G1329gat));
  XOR2_X1   g487(.A(KEYINPUT106), .B(G43gat), .Z(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n646_), .B2(new_n624_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n409_), .A2(new_n403_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n658_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1330gat));
  AOI21_X1  g493(.A(G50gat), .B1(new_n646_), .B2(new_n384_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n384_), .A2(G50gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n658_), .B2(new_n696_), .ZN(G1331gat));
  NOR3_X1   g496(.A1(new_n552_), .A2(new_n641_), .A3(new_n595_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n609_), .A2(G57gat), .A3(new_n386_), .A4(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n464_), .B1(new_n644_), .B2(new_n643_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT107), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n701_), .A2(new_n386_), .A3(new_n601_), .A4(new_n596_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703_));
  INV_X1    g502(.A(G57gat), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n702_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n699_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT109), .B(new_n699_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1332gat));
  AND2_X1   g510(.A1(new_n701_), .A2(new_n601_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n596_), .ZN(new_n713_));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n616_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n609_), .A2(new_n698_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G64gat), .B1(new_n716_), .B2(new_n415_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT48), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n713_), .A2(new_n720_), .A3(new_n624_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G71gat), .B1(new_n716_), .B2(new_n409_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1334gat));
  INV_X1    g523(.A(G78gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n713_), .A2(new_n725_), .A3(new_n384_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G78gat), .B1(new_n716_), .B2(new_n420_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT50), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1335gat));
  AND3_X1   g528(.A1(new_n650_), .A2(new_n651_), .A3(new_n595_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n464_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n552_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n385_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n639_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n712_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n386_), .A2(new_n478_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(G1336gat));
  NAND3_X1  g537(.A1(new_n712_), .A2(new_n616_), .A3(new_n735_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n733_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n616_), .A2(G92gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT110), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n739_), .A2(new_n479_), .B1(new_n740_), .B2(new_n742_), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n733_), .B2(new_n409_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n624_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n736_), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g546(.A1(new_n712_), .A2(new_n475_), .A3(new_n384_), .A4(new_n735_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n730_), .A2(new_n384_), .A3(new_n732_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(G106gat), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n749_), .B2(G106gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n754_), .B(new_n756_), .ZN(G1339gat));
  AOI21_X1  g556(.A(new_n470_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(new_n464_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n530_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT55), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n545_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n533_), .A2(new_n763_), .A3(KEYINPUT55), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT55), .B(new_n472_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT113), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n764_), .A3(new_n766_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n470_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n470_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n759_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n456_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n445_), .A2(new_n771_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n455_), .B2(new_n773_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n774_), .A2(new_n425_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n461_), .B2(new_n460_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n546_), .A2(new_n547_), .A3(new_n470_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n758_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n549_), .A2(KEYINPUT114), .A3(new_n776_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n770_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n606_), .A2(new_n607_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT96), .B1(new_n577_), .B2(new_n578_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n784_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n782_), .A2(new_n783_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n783_), .B1(new_n782_), .B2(new_n787_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n541_), .A2(new_n776_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n767_), .A2(new_n470_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n470_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n581_), .B1(new_n796_), .B2(KEYINPUT58), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n768_), .A2(new_n769_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n791_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT114), .B1(new_n549_), .B2(new_n776_), .ZN(new_n802_));
  MUX2_X1   g601(.A(new_n774_), .B(new_n461_), .S(new_n425_), .Z(new_n803_));
  AOI211_X1 g602(.A(new_n779_), .B(new_n803_), .C1(new_n541_), .C2(new_n548_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n608_), .B1(new_n805_), .B2(new_n770_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n801_), .B1(new_n806_), .B2(KEYINPUT57), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n595_), .B1(new_n790_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n596_), .A2(new_n465_), .A3(new_n552_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT54), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n616_), .A2(new_n384_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n409_), .A2(new_n385_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n811_), .A2(KEYINPUT59), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n790_), .B2(new_n807_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n782_), .A2(new_n787_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT115), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n782_), .A2(new_n783_), .A3(new_n787_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n608_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n782_), .A2(new_n823_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n824_), .A2(new_n785_), .B1(new_n800_), .B2(new_n797_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n822_), .A2(KEYINPUT116), .A3(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n818_), .A2(new_n595_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n810_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(KEYINPUT117), .A3(new_n810_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n814_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n833_), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT119), .B1(new_n833_), .B2(KEYINPUT59), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n641_), .B(new_n816_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(G113gat), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n830_), .A2(new_n831_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT118), .A3(new_n832_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n833_), .A2(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n731_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n837_), .A2(new_n844_), .ZN(G1340gat));
  OAI211_X1 g644(.A(new_n601_), .B(new_n816_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G120gat), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT120), .B1(new_n848_), .B2(G120gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(G120gat), .B1(new_n601_), .B2(new_n848_), .ZN(new_n850_));
  MUX2_X1   g649(.A(new_n849_), .B(KEYINPUT120), .S(new_n850_), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n842_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n847_), .A2(new_n852_), .ZN(G1341gat));
  OAI211_X1 g652(.A(new_n603_), .B(new_n816_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G127gat), .ZN(new_n855_));
  INV_X1    g654(.A(G127gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n842_), .A2(new_n856_), .A3(new_n603_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1342gat));
  INV_X1    g657(.A(new_n835_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n833_), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n815_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n582_), .A2(G134gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT121), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n839_), .A2(new_n608_), .A3(new_n841_), .ZN(new_n864_));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n861_), .A2(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1343gat));
  NOR3_X1   g665(.A1(new_n616_), .A2(new_n624_), .A3(new_n385_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n838_), .A2(new_n384_), .A3(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n464_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n219_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n552_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n220_), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n868_), .A2(new_n595_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT61), .B(G155gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n868_), .B2(new_n581_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n823_), .A2(G162gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n868_), .B2(new_n877_), .ZN(G1347gat));
  NAND2_X1  g677(.A1(new_n616_), .A2(new_n416_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT122), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n811_), .A2(new_n384_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n286_), .B1(new_n881_), .B2(new_n731_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT62), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n881_), .B(KEYINPUT123), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT22), .B(G169gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n731_), .A2(new_n886_), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n887_), .B(KEYINPUT124), .Z(new_n888_));
  OAI21_X1  g687(.A(new_n883_), .B1(new_n885_), .B2(new_n888_), .ZN(G1348gat));
  AOI21_X1  g688(.A(G176gat), .B1(new_n884_), .B2(new_n601_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n838_), .A2(new_n420_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n880_), .A2(new_n287_), .A3(new_n552_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1349gat));
  INV_X1    g692(.A(new_n880_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n891_), .A2(new_n603_), .A3(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(G183gat), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n603_), .A2(new_n290_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n895_), .A2(new_n896_), .B1(new_n884_), .B2(new_n897_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n885_), .B2(new_n581_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n823_), .A2(new_n289_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n885_), .B2(new_n900_), .ZN(G1351gat));
  NOR3_X1   g700(.A1(new_n415_), .A2(new_n624_), .A3(new_n386_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n838_), .A2(new_n384_), .A3(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n464_), .ZN(new_n904_));
  INV_X1    g703(.A(G197gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1352gat));
  NOR2_X1   g705(.A1(new_n903_), .A2(new_n552_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n207_), .ZN(G1353gat));
  NAND2_X1  g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n603_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  OAI22_X1  g710(.A1(new_n903_), .A2(new_n910_), .B1(KEYINPUT125), .B2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(KEYINPUT125), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT126), .Z(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n912_), .A2(new_n915_), .ZN(new_n916_));
  OAI221_X1 g715(.A(new_n914_), .B1(KEYINPUT125), .B2(new_n911_), .C1(new_n903_), .C2(new_n910_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1354gat));
  XNOR2_X1  g717(.A(KEYINPUT127), .B(G218gat), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n903_), .A2(new_n581_), .A3(new_n919_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n903_), .A2(new_n823_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n919_), .ZN(G1355gat));
endmodule


