//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT6), .Z(new_n204_));
  INV_X1    g003(.A(G85gat), .ZN(new_n205_));
  INV_X1    g004(.A(G92gat), .ZN(new_n206_));
  NOR3_X1   g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT9), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT10), .B(G99gat), .Z(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G106gat), .Z(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  INV_X1    g014(.A(new_n203_), .ZN(new_n216_));
  AND2_X1   g015(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n203_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT68), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n227_), .B(new_n228_), .C1(new_n229_), .C2(KEYINPUT7), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n231_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n224_), .A2(new_n226_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n212_), .B(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n215_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n212_), .B(KEYINPUT66), .ZN(new_n238_));
  INV_X1    g037(.A(new_n233_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(new_n204_), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n238_), .A2(new_n240_), .A3(KEYINPUT8), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n214_), .B1(new_n237_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G64gat), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT69), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(KEYINPUT69), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT11), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G71gat), .B(G78gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n244_), .A2(new_n250_), .A3(new_n245_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(KEYINPUT11), .A3(new_n248_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n242_), .A2(new_n254_), .A3(KEYINPUT12), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n253_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n239_), .B1(new_n223_), .B2(KEYINPUT68), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n238_), .B1(new_n257_), .B2(new_n226_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n236_), .A2(new_n215_), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n258_), .A2(new_n215_), .B1(new_n240_), .B2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n256_), .B1(new_n260_), .B2(new_n214_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n255_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n256_), .B(new_n214_), .C1(new_n237_), .C2(new_n241_), .ZN(new_n265_));
  INV_X1    g064(.A(G230gat), .ZN(new_n266_));
  INV_X1    g065(.A(G233gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT71), .B1(new_n264_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n265_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n268_), .B1(new_n272_), .B2(new_n261_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n265_), .A2(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n242_), .A2(new_n254_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n262_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .A4(new_n255_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(new_n273_), .A3(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G120gat), .B(G148gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G176gat), .B(G204gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n284_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n271_), .A2(new_n278_), .A3(new_n273_), .A4(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n285_), .A2(KEYINPUT73), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT73), .B1(new_n285_), .B2(new_n287_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n202_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n287_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n285_), .A2(KEYINPUT73), .A3(new_n287_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT13), .A3(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G15gat), .B(G22gat), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  INV_X1    g097(.A(G8gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G8gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G29gat), .B(G36gat), .Z(new_n305_));
  XOR2_X1   g104(.A(G43gat), .B(G50gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT78), .ZN(new_n309_));
  INV_X1    g108(.A(new_n307_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n303_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G229gat), .A2(G233gat), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n307_), .B(KEYINPUT15), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n303_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n309_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT79), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(KEYINPUT79), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G113gat), .B(G141gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT80), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G169gat), .B(G197gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n314_), .A2(new_n318_), .A3(new_n319_), .A4(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n296_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT21), .ZN(new_n330_));
  AND2_X1   g129(.A1(G197gat), .A2(G204gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G197gat), .ZN(new_n334_));
  INV_X1    g133(.A(G204gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G197gat), .A2(G204gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(KEYINPUT21), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT93), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G211gat), .B(G218gat), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n333_), .A2(new_n338_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n333_), .A2(new_n338_), .A3(new_n340_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT93), .B1(new_n338_), .B2(new_n340_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT24), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(G169gat), .B2(G176gat), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n346_), .A2(KEYINPUT96), .ZN(new_n347_));
  INV_X1    g146(.A(G169gat), .ZN(new_n348_));
  INV_X1    g147(.A(G176gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(KEYINPUT96), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  MUX2_X1   g154(.A(KEYINPUT23), .B(new_n353_), .S(new_n355_), .Z(new_n356_));
  NAND3_X1  g155(.A1(new_n345_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT25), .B(G183gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT26), .B(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n352_), .A2(new_n356_), .A3(new_n357_), .A4(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT98), .ZN(new_n362_));
  OR2_X1    g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT83), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT23), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n355_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n354_), .A2(KEYINPUT23), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n363_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT97), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(G169gat), .B2(G176gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n374_), .A2(KEYINPUT82), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n371_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(KEYINPUT82), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(G169gat), .A3(G176gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT97), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n348_), .A2(KEYINPUT22), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(G169gat), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n381_), .A2(new_n383_), .A3(G176gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AND4_X1   g184(.A1(new_n362_), .A2(new_n370_), .A3(new_n380_), .A4(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n355_), .A2(new_n364_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n384_), .B1(new_n388_), .B2(new_n363_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n362_), .B1(new_n389_), .B2(new_n380_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n344_), .B(new_n361_), .C1(new_n386_), .C2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(KEYINPUT19), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT20), .ZN(new_n394_));
  INV_X1    g193(.A(new_n344_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT26), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT81), .B1(new_n396_), .B2(G190gat), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n358_), .B(new_n397_), .C1(new_n359_), .C2(KEYINPUT81), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n377_), .A2(new_n378_), .A3(new_n350_), .A4(KEYINPUT24), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n398_), .A2(new_n388_), .A3(new_n357_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n354_), .A2(new_n364_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(new_n363_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT84), .B1(new_n348_), .B2(KEYINPUT22), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT22), .B(G169gat), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n349_), .B(new_n403_), .C1(new_n404_), .C2(KEYINPUT84), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n373_), .A2(new_n375_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n394_), .B1(new_n395_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n391_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT99), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT99), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n391_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n361_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n395_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n344_), .A2(new_n407_), .A3(new_n400_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT20), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT95), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n420_), .A3(KEYINPUT20), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n416_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n393_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT18), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  NAND3_X1  g227(.A1(new_n414_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT102), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT102), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n414_), .A2(new_n424_), .A3(new_n431_), .A4(new_n428_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n361_), .A2(new_n344_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n380_), .B2(new_n389_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n395_), .A2(new_n408_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n423_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n428_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n433_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n430_), .A2(new_n432_), .A3(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n414_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n428_), .B1(new_n414_), .B2(new_n424_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n433_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT103), .ZN(new_n447_));
  INV_X1    g246(.A(new_n421_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n420_), .B1(new_n417_), .B2(KEYINPUT20), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n393_), .B1(new_n450_), .B2(new_n416_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n391_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n412_), .B1(new_n391_), .B2(new_n409_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n441_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n429_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT103), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n433_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n443_), .B1(new_n447_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n408_), .B(KEYINPUT30), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G227gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT85), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G43gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G71gat), .B(G99gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n462_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n460_), .A2(new_n461_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n470_), .A3(new_n468_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G127gat), .B(G134gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G113gat), .B(G120gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT87), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n473_), .B(new_n475_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n478_), .B2(KEYINPUT87), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT31), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n472_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(KEYINPUT88), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n469_), .A2(new_n482_), .A3(new_n471_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n483_), .A2(new_n484_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G155gat), .ZN(new_n489_));
  INV_X1    g288(.A(G162gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT90), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(G155gat), .B2(G162gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G155gat), .A2(G162gat), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n491_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT3), .ZN(new_n499_));
  INV_X1    g298(.A(G141gat), .ZN(new_n500_));
  INV_X1    g299(.A(G148gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n495_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n494_), .A2(KEYINPUT1), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT1), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(G155gat), .A3(G162gat), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n507_), .A2(new_n491_), .A3(new_n493_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n500_), .A2(new_n501_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G141gat), .A2(G148gat), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n506_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n479_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n506_), .A2(new_n478_), .A3(new_n514_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(KEYINPUT4), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G225gat), .A2(G233gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT4), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n479_), .A2(new_n521_), .A3(new_n515_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n516_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G1gat), .B(G29gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G85gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT0), .B(G57gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n516_), .A2(KEYINPUT4), .A3(new_n517_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n522_), .A2(new_n520_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n524_), .B(new_n529_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT94), .B(G106gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n496_), .B(KEYINPUT91), .ZN(new_n539_));
  INV_X1    g338(.A(new_n505_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n541_), .A2(new_n495_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n395_), .B(KEYINPUT92), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(new_n545_), .A3(new_n543_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n506_), .A2(new_n543_), .A3(new_n514_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT28), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G22gat), .B(G50gat), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n546_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n544_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n546_), .A2(new_n548_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n544_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n546_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G228gat), .A2(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(G78gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n553_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n538_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n551_), .A2(new_n552_), .A3(new_n544_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n556_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n561_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n553_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n537_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n459_), .A2(new_n488_), .A3(new_n536_), .A4(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n518_), .A2(new_n519_), .A3(new_n522_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n516_), .A2(new_n517_), .A3(new_n520_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n575_), .A2(new_n530_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n534_), .A2(new_n573_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n523_), .A2(KEYINPUT33), .A3(new_n524_), .A4(new_n529_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT100), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n578_), .A2(new_n579_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n581_), .A2(new_n429_), .A3(new_n455_), .A4(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n440_), .A2(KEYINPUT32), .A3(new_n428_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n428_), .A2(KEYINPUT32), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n414_), .A2(new_n424_), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n586_), .A3(new_n535_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n583_), .A2(new_n587_), .B1(new_n570_), .B2(new_n565_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n565_), .A2(new_n536_), .A3(new_n570_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n459_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n572_), .B1(new_n590_), .B2(new_n488_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n242_), .A2(new_n315_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n592_), .B(new_n597_), .C1(new_n310_), .C2(new_n242_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n595_), .A2(new_n596_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT75), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n598_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT36), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n601_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(KEYINPUT37), .A3(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n303_), .B(new_n615_), .Z(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n256_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT76), .Z(new_n618_));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT16), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT17), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT77), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n617_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n622_), .A2(KEYINPUT17), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n623_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n614_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n329_), .A2(new_n591_), .A3(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n633_), .A2(G1gat), .A3(new_n536_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT38), .Z(new_n635_));
  NAND4_X1  g434(.A1(new_n290_), .A2(new_n295_), .A3(new_n328_), .A4(new_n630_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n430_), .A2(new_n432_), .A3(new_n442_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n457_), .B1(new_n456_), .B2(new_n433_), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT103), .B(KEYINPUT27), .C1(new_n455_), .C2(new_n429_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n589_), .B(new_n639_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n582_), .A2(new_n580_), .A3(new_n577_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n456_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n587_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n571_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n488_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n571_), .B(new_n639_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n487_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n649_), .B(new_n536_), .C1(new_n481_), .C2(new_n485_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n606_), .A2(new_n608_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n636_), .A2(new_n637_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n638_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n535_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(KEYINPUT105), .A3(G1gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT105), .B1(new_n657_), .B2(G1gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n635_), .B1(new_n658_), .B2(new_n659_), .ZN(G1324gat));
  OR3_X1    g459(.A1(new_n633_), .A2(G8gat), .A3(new_n459_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  INV_X1    g461(.A(new_n459_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n638_), .A2(new_n654_), .A3(new_n655_), .A4(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G8gat), .B1(new_n664_), .B2(KEYINPUT106), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(KEYINPUT106), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n662_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n667_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n669_), .A2(new_n665_), .A3(KEYINPUT39), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n661_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT40), .B(new_n661_), .C1(new_n668_), .C2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1325gat));
  INV_X1    g474(.A(new_n488_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n633_), .A2(G15gat), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n656_), .A2(new_n488_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(new_n678_), .B2(G15gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(G1326gat));
  XNOR2_X1  g480(.A(new_n571_), .B(KEYINPUT107), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n633_), .A2(G22gat), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n656_), .A2(new_n682_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G22gat), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(KEYINPUT42), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(KEYINPUT42), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1327gat));
  NAND3_X1  g488(.A1(new_n296_), .A2(new_n328_), .A3(new_n629_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n652_), .B2(new_n614_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n692_), .B(new_n613_), .C1(new_n647_), .C2(new_n651_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n690_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT108), .B1(new_n694_), .B2(KEYINPUT44), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n692_), .B1(new_n591_), .B2(new_n613_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n693_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n696_), .B(new_n697_), .C1(new_n700_), .C2(new_n690_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n296_), .A2(new_n328_), .A3(new_n629_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n702_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n691_), .A2(new_n693_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n706_), .A2(KEYINPUT109), .A3(KEYINPUT44), .A4(new_n702_), .ZN(new_n707_));
  AOI22_X1  g506(.A1(new_n695_), .A2(new_n701_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(G29gat), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n536_), .A2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n630_), .A2(new_n609_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT110), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n329_), .A2(new_n712_), .A3(new_n591_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT111), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n329_), .A2(new_n712_), .A3(new_n715_), .A4(new_n591_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(new_n535_), .A3(new_n716_), .ZN(new_n717_));
  AOI22_X1  g516(.A1(new_n708_), .A2(new_n710_), .B1(new_n709_), .B2(new_n717_), .ZN(G1328gat));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  INV_X1    g518(.A(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n708_), .B2(new_n663_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n459_), .A2(G36gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n714_), .A2(new_n716_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n719_), .B1(new_n721_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n701_), .A2(new_n695_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n705_), .A2(new_n707_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n663_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G36gat), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n723_), .B(KEYINPUT45), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(KEYINPUT46), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n726_), .A2(new_n732_), .ZN(G1329gat));
  NAND4_X1  g532(.A1(new_n727_), .A2(new_n728_), .A3(G43gat), .A4(new_n488_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n714_), .A2(new_n488_), .A3(new_n716_), .ZN(new_n735_));
  INV_X1    g534(.A(G43gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT47), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n740_), .A3(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1330gat));
  INV_X1    g541(.A(G50gat), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n571_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n714_), .A2(new_n682_), .A3(new_n716_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n708_), .A2(new_n744_), .B1(new_n743_), .B2(new_n745_), .ZN(G1331gat));
  INV_X1    g545(.A(new_n296_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n632_), .A2(new_n747_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT112), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT112), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n652_), .A2(new_n328_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(G57gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n535_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n296_), .A2(new_n328_), .A3(new_n629_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n654_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n756_), .A2(KEYINPUT113), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(KEYINPUT113), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n535_), .A3(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n759_), .B2(new_n753_), .ZN(G1332gat));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n663_), .A3(new_n758_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(G64gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G64gat), .ZN(new_n764_));
  INV_X1    g563(.A(new_n752_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n459_), .A2(G64gat), .ZN(new_n766_));
  OAI22_X1  g565(.A1(new_n763_), .A2(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(G1333gat));
  NAND3_X1  g566(.A1(new_n757_), .A2(new_n488_), .A3(new_n758_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(G71gat), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G71gat), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n676_), .A2(G71gat), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n770_), .A2(new_n771_), .B1(new_n765_), .B2(new_n772_), .ZN(G1334gat));
  NAND3_X1  g572(.A1(new_n752_), .A2(new_n560_), .A3(new_n682_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n757_), .A2(new_n682_), .A3(new_n758_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(G78gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G78gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1335gat));
  NOR3_X1   g578(.A1(new_n296_), .A2(new_n328_), .A3(new_n630_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n706_), .A2(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n535_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n712_), .A2(new_n747_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n751_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n535_), .A2(new_n205_), .ZN(new_n785_));
  OAI22_X1  g584(.A1(new_n782_), .A2(new_n205_), .B1(new_n784_), .B2(new_n785_), .ZN(G1336gat));
  AND2_X1   g585(.A1(new_n781_), .A2(new_n663_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n663_), .A2(new_n206_), .ZN(new_n788_));
  OAI22_X1  g587(.A1(new_n787_), .A2(new_n206_), .B1(new_n784_), .B2(new_n788_), .ZN(G1337gat));
  INV_X1    g588(.A(new_n209_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n784_), .A2(new_n790_), .A3(new_n676_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n781_), .A2(new_n488_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G99gat), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT116), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(KEYINPUT51), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT115), .B1(new_n793_), .B2(KEYINPUT116), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n793_), .B2(KEYINPUT115), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n796_), .B1(new_n797_), .B2(new_n799_), .ZN(G1338gat));
  INV_X1    g599(.A(new_n571_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n783_), .A2(new_n210_), .A3(new_n801_), .A4(new_n751_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n781_), .A2(new_n801_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(G106gat), .ZN(new_n805_));
  AOI211_X1 g604(.A(KEYINPUT52), .B(new_n228_), .C1(new_n781_), .C2(new_n801_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT53), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(new_n802_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1339gat));
  XOR2_X1   g610(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n812_));
  NAND2_X1  g611(.A1(new_n328_), .A2(new_n287_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n264_), .A2(new_n270_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n276_), .A2(new_n265_), .A3(new_n255_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n814_), .A2(KEYINPUT55), .B1(new_n268_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n271_), .A2(new_n817_), .A3(new_n278_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n284_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n284_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n813_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n313_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n309_), .A2(new_n825_), .A3(new_n316_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n325_), .B(new_n826_), .C1(new_n312_), .C2(new_n825_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n327_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT118), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n828_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n824_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n812_), .B1(new_n833_), .B2(new_n653_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n824_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n293_), .A2(new_n294_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n831_), .B1(new_n836_), .B2(new_n828_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n832_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n835_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n609_), .A2(KEYINPUT57), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT120), .B1(new_n833_), .B2(new_n841_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n822_), .A2(new_n823_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n828_), .A2(new_n287_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n614_), .B1(new_n847_), .B2(KEYINPUT58), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n846_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n834_), .A2(new_n843_), .A3(new_n844_), .A4(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n629_), .A2(new_n328_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n290_), .A2(new_n295_), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n290_), .A2(new_n295_), .A3(KEYINPUT117), .A4(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n614_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT54), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n862_), .A3(new_n614_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n853_), .A2(new_n629_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n488_), .A2(new_n535_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n648_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT59), .B1(new_n864_), .B2(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n866_), .A2(KEYINPUT121), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n866_), .A2(KEYINPUT121), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n869_), .A2(new_n870_), .A3(KEYINPUT59), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n843_), .A2(new_n844_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n839_), .A2(new_n609_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n873_), .A2(new_n812_), .B1(new_n848_), .B2(new_n851_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n630_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n861_), .A2(new_n863_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n871_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n868_), .A2(new_n328_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G113gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n853_), .A2(new_n629_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n861_), .A2(new_n863_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n866_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n328_), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n883_), .A2(G113gat), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n879_), .A2(new_n885_), .ZN(G1340gat));
  NAND3_X1  g685(.A1(new_n868_), .A2(new_n747_), .A3(new_n877_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G120gat), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n296_), .A2(KEYINPUT60), .ZN(new_n889_));
  MUX2_X1   g688(.A(new_n889_), .B(KEYINPUT60), .S(G120gat), .Z(new_n890_));
  NAND3_X1  g689(.A1(new_n882_), .A2(new_n866_), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n864_), .A2(new_n867_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(KEYINPUT122), .A3(new_n890_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n888_), .A2(new_n896_), .ZN(G1341gat));
  NAND3_X1  g696(.A1(new_n868_), .A2(new_n630_), .A3(new_n877_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G127gat), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n883_), .A2(G127gat), .A3(new_n629_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1342gat));
  AOI21_X1  g700(.A(G134gat), .B1(new_n894_), .B2(new_n653_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n868_), .A2(new_n877_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT123), .B(G134gat), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n614_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n903_), .B2(new_n905_), .ZN(G1343gat));
  NAND4_X1  g705(.A1(new_n676_), .A2(new_n535_), .A3(new_n801_), .A4(new_n459_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n882_), .A2(new_n328_), .A3(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g709(.A1(new_n864_), .A2(new_n907_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT124), .B(G148gat), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n911_), .A2(new_n747_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n911_), .B2(new_n747_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1345gat));
  NAND3_X1  g714(.A1(new_n882_), .A2(new_n630_), .A3(new_n908_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT61), .B(G155gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  NAND3_X1  g717(.A1(new_n911_), .A2(new_n490_), .A3(new_n653_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n864_), .A2(new_n614_), .A3(new_n907_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n490_), .B2(new_n920_), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n459_), .A2(new_n650_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n682_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI211_X1 g726(.A(KEYINPUT62), .B(G169gat), .C1(new_n927_), .C2(new_n884_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n864_), .A2(new_n884_), .A3(new_n925_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n348_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n404_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(new_n931_), .A3(new_n932_), .ZN(G1348gat));
  AOI21_X1  g732(.A(G176gat), .B1(new_n926_), .B2(new_n747_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n864_), .A2(new_n801_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n296_), .A2(new_n923_), .A3(new_n349_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n934_), .B1(new_n935_), .B2(new_n936_), .ZN(G1349gat));
  NOR2_X1   g736(.A1(new_n923_), .A2(new_n629_), .ZN(new_n938_));
  AOI21_X1  g737(.A(G183gat), .B1(new_n935_), .B2(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n629_), .A2(new_n358_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n926_), .B2(new_n940_), .ZN(G1350gat));
  NAND2_X1  g740(.A1(new_n653_), .A2(new_n359_), .ZN(new_n942_));
  XOR2_X1   g741(.A(new_n942_), .B(KEYINPUT126), .Z(new_n943_));
  NAND2_X1  g742(.A1(new_n926_), .A2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  INV_X1    g744(.A(G190gat), .ZN(new_n946_));
  AOI211_X1 g745(.A(new_n945_), .B(new_n946_), .C1(new_n926_), .C2(new_n613_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n613_), .B(new_n924_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n948_));
  AOI21_X1  g747(.A(KEYINPUT125), .B1(new_n948_), .B2(G190gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n944_), .B1(new_n947_), .B2(new_n949_), .ZN(G1351gat));
  NAND3_X1  g749(.A1(new_n663_), .A2(new_n676_), .A3(new_n589_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n882_), .A2(G197gat), .A3(new_n328_), .A4(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n864_), .A2(new_n951_), .ZN(new_n956_));
  NAND4_X1  g755(.A1(new_n956_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n328_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n882_), .A2(new_n328_), .A3(new_n952_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n334_), .ZN(new_n959_));
  AND3_X1   g758(.A1(new_n955_), .A2(new_n957_), .A3(new_n959_), .ZN(G1352gat));
  INV_X1    g759(.A(new_n956_), .ZN(new_n961_));
  OAI21_X1  g760(.A(G204gat), .B1(new_n961_), .B2(new_n296_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n956_), .A2(new_n335_), .A3(new_n747_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1353gat));
  OR2_X1    g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(new_n956_), .B2(new_n630_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n961_), .A2(new_n629_), .ZN(new_n967_));
  XOR2_X1   g766(.A(KEYINPUT63), .B(G211gat), .Z(new_n968_));
  AOI21_X1  g767(.A(new_n966_), .B1(new_n967_), .B2(new_n968_), .ZN(G1354gat));
  OAI21_X1  g768(.A(G218gat), .B1(new_n961_), .B2(new_n614_), .ZN(new_n970_));
  INV_X1    g769(.A(G218gat), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n956_), .A2(new_n971_), .A3(new_n653_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n970_), .A2(new_n972_), .ZN(G1355gat));
endmodule


