//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT17), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G155gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT16), .ZN(new_n205_));
  XOR2_X1   g004(.A(G183gat), .B(G211gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT79), .B(G8gat), .Z(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(new_n209_), .B2(new_n202_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n208_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n211_), .A3(new_n208_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(G231gat), .A2(G233gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G57gat), .B(G64gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT11), .ZN(new_n219_));
  XOR2_X1   g018(.A(G71gat), .B(G78gat), .Z(new_n220_));
  OR2_X1    g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n218_), .A2(KEYINPUT11), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n220_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  AOI211_X1 g025(.A(new_n203_), .B(new_n207_), .C1(new_n217_), .C2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(new_n226_), .B2(new_n217_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n207_), .B(new_n203_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n217_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n230_), .B2(new_n224_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(new_n224_), .B2(new_n230_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT12), .ZN(new_n235_));
  INV_X1    g034(.A(G85gat), .ZN(new_n236_));
  INV_X1    g035(.A(G92gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G85gat), .A2(G92gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n238_), .B(new_n239_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G99gat), .A2(G106gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT6), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT6), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G99gat), .A3(G106gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT7), .ZN(new_n249_));
  INV_X1    g048(.A(G99gat), .ZN(new_n250_));
  INV_X1    g049(.A(G106gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n247_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n242_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n247_), .A2(KEYINPUT65), .A3(new_n248_), .A4(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n238_), .A2(new_n239_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n244_), .A2(new_n246_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n248_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n255_), .A2(new_n256_), .B1(KEYINPUT8), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT9), .ZN(new_n263_));
  INV_X1    g062(.A(new_n239_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n238_), .B(new_n263_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n238_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n239_), .ZN(new_n267_));
  OR2_X1    g066(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n251_), .A3(new_n269_), .ZN(new_n270_));
  AND4_X1   g069(.A1(new_n247_), .A2(new_n266_), .A3(new_n267_), .A4(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n262_), .A2(new_n271_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n226_), .A2(new_n235_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n262_), .B2(new_n271_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n254_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n242_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n256_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n261_), .A2(KEYINPUT8), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n271_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(KEYINPUT67), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(new_n224_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G230gat), .ZN(new_n285_));
  INV_X1    g084(.A(G233gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n224_), .B1(new_n276_), .B2(new_n283_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT12), .ZN(new_n293_));
  INV_X1    g092(.A(new_n224_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT67), .B1(new_n281_), .B2(new_n282_), .ZN(new_n295_));
  AOI211_X1 g094(.A(new_n275_), .B(new_n271_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT69), .B1(new_n297_), .B2(new_n235_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n274_), .B(new_n290_), .C1(new_n293_), .C2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n284_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n287_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n292_), .B1(new_n291_), .B2(KEYINPUT12), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n297_), .A2(KEYINPUT69), .A3(new_n235_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n273_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(KEYINPUT70), .A3(new_n290_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n301_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G176gat), .B(G204gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT72), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G120gat), .B(G148gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n314_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n301_), .A2(new_n307_), .A3(new_n303_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT13), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT84), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G113gat), .B(G141gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT82), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G169gat), .B(G197gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G229gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT80), .ZN(new_n330_));
  INV_X1    g129(.A(new_n214_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(new_n212_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G29gat), .B(G36gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G43gat), .B(G50gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n330_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n215_), .A2(KEYINPUT80), .A3(new_n335_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n335_), .B(KEYINPUT15), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n332_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n329_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n331_), .A2(new_n212_), .A3(new_n335_), .ZN(new_n343_));
  AOI211_X1 g142(.A(new_n328_), .B(new_n343_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n327_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n326_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n342_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n327_), .B1(new_n325_), .B2(KEYINPUT83), .ZN(new_n349_));
  INV_X1    g148(.A(new_n343_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n339_), .A2(new_n329_), .A3(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n321_), .B1(new_n347_), .B2(new_n353_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n337_), .A2(new_n338_), .B1(new_n332_), .B2(new_n340_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n351_), .B1(new_n329_), .B2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT83), .B1(new_n356_), .B2(new_n327_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT84), .B(new_n352_), .C1(new_n357_), .C2(new_n326_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n320_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G190gat), .B(G218gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G134gat), .B(G162gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT36), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT76), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT35), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n368_));
  NAND2_X1  g167(.A1(G232gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT15), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n335_), .B(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT74), .B1(new_n272_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n340_), .B(new_n374_), .C1(new_n262_), .C2(new_n271_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n276_), .A2(new_n335_), .A3(new_n283_), .ZN(new_n377_));
  AOI211_X1 g176(.A(new_n367_), .B(new_n370_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n370_), .A2(new_n367_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n370_), .A2(new_n367_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n376_), .A2(new_n380_), .A3(new_n381_), .A4(new_n377_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n366_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n376_), .A2(new_n381_), .A3(new_n377_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n379_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n364_), .A2(KEYINPUT36), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n382_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(G85gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(G155gat), .A2(G162gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n399_), .B(KEYINPUT3), .Z(new_n400_));
  NAND2_X1  g199(.A1(G141gat), .A2(G148gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n401_), .B(KEYINPUT2), .Z(new_n402_));
  OAI211_X1 g201(.A(new_n397_), .B(new_n398_), .C1(new_n400_), .C2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT1), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n398_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n397_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n399_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n401_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G127gat), .B(G134gat), .Z(new_n411_));
  XOR2_X1   g210(.A(G113gat), .B(G120gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(KEYINPUT4), .A3(new_n416_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT99), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n418_), .B1(new_n415_), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n421_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n394_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n420_), .A2(new_n423_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT99), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n429_), .A2(new_n393_), .A3(new_n419_), .A4(new_n424_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT89), .ZN(new_n432_));
  XOR2_X1   g231(.A(G71gat), .B(G99gat), .Z(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G43gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(G15gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n434_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G183gat), .A2(G190gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT23), .ZN(new_n441_));
  OR3_X1    g240(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(KEYINPUT86), .A2(G190gat), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n444_), .A2(KEYINPUT26), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(KEYINPUT26), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT25), .B1(KEYINPUT85), .B2(G183gat), .ZN(new_n447_));
  AND3_X1   g246(.A1(KEYINPUT85), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n445_), .B(new_n446_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G169gat), .A2(G176gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n443_), .B(new_n449_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT22), .B(G169gat), .Z(new_n455_));
  OR2_X1    g254(.A1(new_n455_), .A2(G176gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n441_), .B1(G183gat), .B2(G190gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n450_), .B(KEYINPUT87), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT30), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n454_), .A2(KEYINPUT30), .A3(new_n459_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n439_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n439_), .A3(new_n463_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n438_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n438_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT31), .B1(new_n467_), .B2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n468_), .B2(new_n464_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT31), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n472_), .B(new_n473_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n432_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n413_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n471_), .A2(new_n474_), .A3(new_n432_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n413_), .B1(new_n480_), .B2(new_n475_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n431_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G197gat), .B(G204gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT21), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G211gat), .B(G218gat), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n485_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n489_), .A3(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n410_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT91), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n483_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G228gat), .A2(G233gat), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n488_), .A2(new_n490_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n497_), .B1(new_n409_), .B2(KEYINPUT29), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n498_), .B2(KEYINPUT92), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n483_), .B(new_n496_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G78gat), .B(G106gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n500_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n409_), .A2(KEYINPUT29), .ZN(new_n508_));
  XOR2_X1   g307(.A(G22gat), .B(G50gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT28), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n508_), .B(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n503_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n511_), .B1(new_n512_), .B2(KEYINPUT93), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n505_), .A2(KEYINPUT93), .A3(new_n506_), .A4(new_n511_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n452_), .A2(KEYINPUT97), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT97), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n458_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n456_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n520_), .B2(new_n456_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n457_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT25), .B(G183gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(G190gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n453_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n525_), .A2(new_n526_), .B1(new_n527_), .B2(new_n450_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n443_), .A2(KEYINPUT95), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n441_), .A2(new_n442_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT95), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n528_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT96), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n530_), .B(new_n531_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT96), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n528_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n524_), .A2(new_n534_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n491_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT20), .B1(new_n460_), .B2(new_n491_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G226gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G8gat), .B(G36gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT18), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G64gat), .B(G92gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(KEYINPUT20), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n551_), .B1(new_n460_), .B2(new_n491_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n545_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n524_), .A2(new_n534_), .A3(new_n497_), .A4(new_n537_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n546_), .A2(KEYINPUT103), .A3(new_n550_), .A4(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n540_), .B1(new_n538_), .B2(new_n491_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n556_), .B(new_n550_), .C1(new_n558_), .C2(new_n553_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT103), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  AOI211_X1 g361(.A(new_n540_), .B(new_n545_), .C1(new_n538_), .C2(new_n491_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n524_), .A2(new_n497_), .A3(new_n533_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n553_), .B1(new_n564_), .B2(new_n552_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT102), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n558_), .A2(new_n553_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT102), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n550_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT27), .B1(new_n562_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n556_), .B1(new_n558_), .B2(new_n553_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n550_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n559_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT27), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n516_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n482_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n571_), .A2(new_n577_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n431_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n572_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n550_), .A2(KEYINPUT32), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n431_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n583_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(KEYINPUT100), .A2(KEYINPUT33), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n430_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n419_), .A2(new_n424_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n587_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n589_), .A2(new_n393_), .A3(new_n429_), .A4(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n418_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n393_), .B1(new_n417_), .B2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n415_), .B2(new_n422_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n420_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n595_), .A2(KEYINPUT101), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(KEYINPUT101), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n591_), .A3(new_n598_), .ZN(new_n599_));
  OAI22_X1  g398(.A1(new_n585_), .A2(new_n586_), .B1(new_n599_), .B2(new_n575_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n516_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n580_), .A2(new_n581_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n479_), .A2(new_n481_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n579_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  AND4_X1   g403(.A1(new_n234_), .A2(new_n361_), .A3(new_n389_), .A4(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n202_), .B1(new_n605_), .B2(new_n431_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT77), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n384_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n388_), .A2(KEYINPUT75), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT75), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n386_), .A2(new_n610_), .A3(new_n387_), .A4(new_n382_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT77), .B(new_n366_), .C1(new_n378_), .C2(new_n383_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n608_), .A2(new_n609_), .A3(new_n611_), .A4(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT37), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n384_), .A2(new_n615_), .A3(new_n388_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT78), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT78), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n384_), .A2(new_n618_), .A3(new_n615_), .A4(new_n388_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(new_n233_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n361_), .A2(new_n623_), .A3(new_n604_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT104), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT104), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n361_), .A2(new_n626_), .A3(new_n604_), .A4(new_n623_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n431_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(G1gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n606_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n625_), .A2(KEYINPUT38), .A3(new_n627_), .A4(new_n629_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(new_n634_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1324gat));
  INV_X1    g438(.A(new_n565_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n568_), .B1(new_n567_), .B2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n563_), .A2(KEYINPUT102), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n573_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n561_), .A3(new_n557_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n576_), .B1(new_n644_), .B2(KEYINPUT27), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n625_), .A2(new_n209_), .A3(new_n645_), .A4(new_n627_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n389_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n516_), .A2(new_n628_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n588_), .A2(new_n591_), .A3(new_n598_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n575_), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n430_), .A2(new_n427_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT32), .B(new_n550_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n649_), .A2(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  OAI22_X1  g452(.A1(new_n645_), .A2(new_n648_), .B1(new_n653_), .B2(new_n516_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n603_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n647_), .B1(new_n656_), .B2(new_n579_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n657_), .A2(new_n234_), .A3(new_n361_), .A4(new_n645_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G8gat), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT107), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(new_n662_), .A3(G8gat), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n661_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n646_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT40), .B(new_n646_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1325gat));
  NAND2_X1  g469(.A1(new_n605_), .A2(new_n603_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n671_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT41), .B1(new_n671_), .B2(G15gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n625_), .A2(new_n627_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n603_), .A2(new_n436_), .ZN(new_n675_));
  OAI22_X1  g474(.A1(new_n672_), .A2(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n605_), .A2(new_n516_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G22gat), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n601_), .A2(G22gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n674_), .B2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n389_), .A2(new_n234_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n361_), .A2(new_n604_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(G29gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n431_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n361_), .A2(new_n233_), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n654_), .A2(new_n655_), .B1(new_n578_), .B2(new_n482_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n693_), .B2(new_n621_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n604_), .A2(new_n695_), .A3(new_n622_), .ZN(new_n696_));
  AOI211_X1 g495(.A(new_n691_), .B(new_n692_), .C1(new_n694_), .C2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n694_), .A2(new_n696_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n692_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT44), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n431_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n690_), .B1(new_n702_), .B2(G29gat), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT110), .B(new_n688_), .C1(new_n701_), .C2(new_n431_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n689_), .B1(new_n703_), .B2(new_n704_), .ZN(G1328gat));
  NAND2_X1  g504(.A1(new_n698_), .A2(new_n699_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n691_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n698_), .A2(KEYINPUT44), .A3(new_n699_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n645_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G36gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n580_), .A2(G36gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n687_), .A2(KEYINPUT112), .A3(new_n711_), .ZN(new_n712_));
  XOR2_X1   g511(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n713_));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n714_));
  INV_X1    g513(.A(new_n711_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n686_), .B2(new_n715_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n712_), .A2(new_n713_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n713_), .B1(new_n712_), .B2(new_n716_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n710_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n710_), .B2(new_n719_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  AOI21_X1  g522(.A(G43gat), .B1(new_n687_), .B2(new_n603_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n603_), .A2(G43gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n701_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n687_), .B2(new_n516_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n516_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n701_), .B2(new_n730_), .ZN(G1331gat));
  XNOR2_X1  g530(.A(new_n318_), .B(KEYINPUT13), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n693_), .A2(new_n359_), .A3(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n623_), .ZN(new_n734_));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n431_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n732_), .A2(new_n359_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n657_), .A2(new_n234_), .A3(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(new_n431_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n736_), .B1(new_n739_), .B2(new_n735_), .ZN(G1332gat));
  INV_X1    g539(.A(G64gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n738_), .B2(new_n645_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n734_), .A2(new_n741_), .A3(new_n645_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n738_), .B2(new_n603_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT49), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n734_), .A2(new_n747_), .A3(new_n603_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n738_), .B2(new_n516_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n734_), .A2(new_n752_), .A3(new_n516_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1335gat));
  NOR3_X1   g556(.A1(new_n693_), .A2(KEYINPUT43), .A3(new_n621_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n695_), .B1(new_n604_), .B2(new_n622_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT116), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n737_), .A2(new_n233_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n694_), .A2(new_n763_), .A3(new_n696_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n628_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n733_), .A2(new_n685_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n236_), .A3(new_n431_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1336gat));
  OAI21_X1  g568(.A(G92gat), .B1(new_n765_), .B2(new_n580_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n237_), .A3(new_n645_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1337gat));
  NAND4_X1  g571(.A1(new_n760_), .A2(new_n603_), .A3(new_n762_), .A4(new_n764_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G99gat), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n603_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n733_), .A2(new_n685_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT117), .B1(new_n778_), .B2(KEYINPUT51), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n776_), .B1(new_n773_), .B2(G99gat), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n785_));
  AND4_X1   g584(.A1(new_n784_), .A2(new_n774_), .A3(new_n777_), .A4(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n780_), .B2(new_n785_), .ZN(new_n787_));
  OAI22_X1  g586(.A1(new_n779_), .A2(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n767_), .A2(new_n251_), .A3(new_n516_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n761_), .A2(new_n601_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n698_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n792_), .B2(G106gat), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT52), .B(new_n251_), .C1(new_n698_), .C2(new_n791_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n789_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI211_X1 g595(.A(new_n233_), .B(new_n359_), .C1(new_n614_), .C2(new_n620_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n732_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(new_n732_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n359_), .A2(new_n317_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n301_), .A2(new_n803_), .A3(new_n307_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n273_), .B(new_n289_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n284_), .B(new_n274_), .C1(new_n293_), .C2(new_n298_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n805_), .A2(KEYINPUT55), .B1(new_n806_), .B2(new_n287_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n314_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n314_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n802_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n355_), .A2(new_n328_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n339_), .A2(new_n328_), .A3(new_n350_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n326_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n326_), .B2(new_n356_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n318_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n389_), .B1(new_n813_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n359_), .A2(new_n317_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n314_), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n810_), .B(new_n316_), .C1(new_n804_), .C2(new_n807_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n647_), .B1(new_n826_), .B2(new_n818_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT57), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n317_), .A2(new_n817_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n621_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT58), .B(new_n830_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n822_), .A2(new_n828_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n801_), .B1(new_n836_), .B2(new_n233_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n578_), .A2(new_n603_), .A3(new_n431_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(G113gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n359_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n838_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n820_), .A2(new_n821_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n234_), .B1(new_n845_), .B2(new_n828_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT59), .B(new_n844_), .C1(new_n846_), .C2(new_n801_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n360_), .B1(new_n843_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n841_), .B1(new_n848_), .B2(new_n840_), .ZN(G1340gat));
  AOI21_X1  g648(.A(new_n732_), .B1(new_n843_), .B2(new_n847_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT120), .B(G120gat), .Z(new_n851_));
  AOI21_X1  g650(.A(new_n829_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n622_), .B1(new_n852_), .B2(KEYINPUT58), .ZN(new_n853_));
  INV_X1    g652(.A(new_n834_), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n853_), .A2(new_n854_), .B1(new_n827_), .B2(KEYINPUT57), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n820_), .A2(new_n821_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n233_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n801_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n844_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n851_), .B1(new_n732_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(KEYINPUT60), .B2(new_n851_), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n850_), .A2(new_n851_), .B1(new_n860_), .B2(new_n862_), .ZN(G1341gat));
  NAND2_X1  g662(.A1(new_n234_), .A2(G127gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT121), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT59), .B1(new_n859_), .B2(new_n844_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n837_), .A2(new_n842_), .A3(new_n838_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(G127gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n860_), .B2(new_n233_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(KEYINPUT122), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872_));
  INV_X1    g671(.A(new_n865_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n843_), .B2(new_n847_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G127gat), .B1(new_n839_), .B2(new_n234_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n871_), .A2(new_n876_), .ZN(G1342gat));
  INV_X1    g676(.A(G134gat), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n878_), .B(new_n621_), .C1(new_n843_), .C2(new_n847_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n860_), .B2(new_n389_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT123), .B(new_n878_), .C1(new_n860_), .C2(new_n389_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n882_), .B2(new_n883_), .ZN(G1343gat));
  NAND4_X1  g683(.A1(new_n655_), .A2(new_n516_), .A3(new_n580_), .A4(new_n431_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n837_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n359_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n320_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n234_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n886_), .B2(new_n647_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n622_), .A2(G162gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT124), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n886_), .B2(new_n896_), .ZN(G1347gat));
  AND2_X1   g696(.A1(new_n482_), .A2(new_n645_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n359_), .ZN(new_n899_));
  XOR2_X1   g698(.A(new_n899_), .B(KEYINPUT125), .Z(new_n900_));
  NAND3_X1  g699(.A1(new_n859_), .A2(new_n601_), .A3(new_n900_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n902_));
  AND3_X1   g701(.A1(new_n901_), .A2(G169gat), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n901_), .B2(G169gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n859_), .A2(new_n601_), .A3(new_n898_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n360_), .A2(new_n455_), .ZN(new_n906_));
  OAI22_X1  g705(.A1(new_n903_), .A2(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1348gat));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n732_), .ZN(new_n908_));
  INV_X1    g707(.A(G176gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1349gat));
  NOR2_X1   g709(.A1(new_n905_), .A2(new_n233_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(G183gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n905_), .A2(new_n233_), .A3(new_n525_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n905_), .B2(new_n621_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n647_), .A2(new_n526_), .ZN(new_n916_));
  XOR2_X1   g715(.A(new_n916_), .B(KEYINPUT127), .Z(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n905_), .B2(new_n917_), .ZN(G1351gat));
  NAND4_X1  g717(.A1(new_n655_), .A2(new_n516_), .A3(new_n645_), .A4(new_n628_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n837_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n359_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n320_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g723(.A(KEYINPUT63), .B(G211gat), .C1(new_n920_), .C2(new_n234_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n837_), .A2(new_n233_), .A3(new_n919_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT63), .B(G211gat), .Z(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(G1354gat));
  INV_X1    g727(.A(G218gat), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n920_), .A2(new_n929_), .A3(new_n647_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n837_), .A2(new_n621_), .A3(new_n919_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n929_), .ZN(G1355gat));
endmodule


