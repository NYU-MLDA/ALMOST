//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT86), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT86), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n209_), .A3(KEYINPUT23), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT93), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n207_), .A2(new_n209_), .A3(KEYINPUT93), .A4(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n206_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT91), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT91), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G169gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT88), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G169gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n226_), .B1(KEYINPUT22), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT22), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT89), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT89), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT22), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n227_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT90), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT89), .B(KEYINPUT22), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n240_), .A2(KEYINPUT90), .A3(new_n227_), .ZN(new_n241_));
  OAI211_X1 g040(.A(KEYINPUT92), .B(new_n232_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n238_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT90), .B1(new_n240_), .B2(new_n227_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT92), .B1(new_n246_), .B2(new_n232_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n220_), .B(new_n221_), .C1(new_n243_), .C2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n207_), .A2(new_n209_), .A3(new_n216_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n215_), .A2(KEYINPUT23), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT24), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n227_), .A3(new_n222_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT87), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT87), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT25), .B(G183gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G190gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n252_), .B1(G169gat), .B2(G176gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n227_), .A2(new_n222_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n258_), .A2(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n255_), .A2(new_n257_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n248_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT30), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G71gat), .B(G99gat), .ZN(new_n266_));
  INV_X1    g065(.A(G43gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G227gat), .A2(G233gat), .ZN(new_n269_));
  INV_X1    g068(.A(G15gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n268_), .B(new_n271_), .Z(new_n272_));
  OR2_X1    g071(.A1(new_n265_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT31), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(new_n272_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n274_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n205_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(new_n276_), .A3(new_n204_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G8gat), .B(G36gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT18), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G64gat), .B(G92gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT20), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT98), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n294_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT99), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n298_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT99), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n295_), .A4(new_n296_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n292_), .A2(new_n296_), .A3(new_n294_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n248_), .A2(new_n263_), .A3(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n218_), .A2(new_n253_), .A3(new_n262_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n251_), .A2(new_n219_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n226_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n221_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n304_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI211_X1 g115(.A(new_n288_), .B(new_n291_), .C1(new_n307_), .C2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n291_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n248_), .A2(new_n263_), .A3(new_n315_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n288_), .B1(new_n314_), .B2(new_n306_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n287_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n307_), .A2(new_n316_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(KEYINPUT20), .A3(new_n318_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n320_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n291_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n326_), .A3(new_n286_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT107), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G22gat), .B(G50gat), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  AND3_X1   g134(.A1(KEYINPUT95), .A2(G155gat), .A3(G162gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT95), .B1(G155gat), .B2(G162gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT1), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT95), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n342_));
  NAND3_X1  g141(.A1(KEYINPUT95), .A2(G155gat), .A3(G162gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G155gat), .ZN(new_n345_));
  INV_X1    g144(.A(G162gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n338_), .A2(new_n344_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT94), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT94), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(G141gat), .ZN(new_n353_));
  INV_X1    g152(.A(G148gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n350_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n348_), .A2(new_n356_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n341_), .A2(new_n343_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT96), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT96), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n361_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n360_), .A2(new_n362_), .A3(new_n363_), .A4(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n350_), .A2(new_n352_), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n358_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n335_), .B1(new_n357_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G233gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(KEYINPUT97), .A2(G228gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(KEYINPUT97), .A2(G228gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n372_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n306_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n315_), .B2(new_n370_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n334_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n357_), .A2(new_n369_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(KEYINPUT29), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT28), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n378_), .A2(new_n379_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n380_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n390_), .A2(new_n382_), .A3(new_n333_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n385_), .A2(new_n388_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n388_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n328_), .A2(KEYINPUT107), .A3(new_n329_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n323_), .A2(KEYINPUT20), .A3(new_n291_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n325_), .A2(new_n318_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT106), .B1(new_n398_), .B2(new_n286_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT106), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n396_), .A2(new_n397_), .A3(new_n400_), .A4(new_n287_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n399_), .A2(KEYINPUT27), .A3(new_n327_), .A4(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n332_), .A2(new_n394_), .A3(new_n395_), .A4(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n386_), .A2(new_n205_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n357_), .A2(new_n369_), .A3(new_n204_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(KEYINPUT4), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n204_), .B1(new_n357_), .B2(new_n369_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n357_), .A2(new_n369_), .A3(new_n204_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n412_), .A2(new_n408_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n407_), .ZN(new_n414_));
  INV_X1    g213(.A(G85gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT0), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n416_), .A2(KEYINPUT0), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n418_), .A2(G57gat), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G57gat), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n416_), .A2(KEYINPUT0), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n417_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n415_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(G57gat), .B1(new_n418_), .B2(new_n419_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n422_), .A2(new_n421_), .A3(new_n417_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(G85gat), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n411_), .A2(new_n414_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT104), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n411_), .A2(new_n414_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(new_n427_), .A3(new_n424_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n411_), .A2(new_n414_), .A3(KEYINPUT104), .A4(new_n428_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n282_), .A2(new_n403_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n435_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n398_), .A2(KEYINPUT32), .A3(new_n286_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n286_), .A2(KEYINPUT32), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT103), .ZN(new_n442_));
  INV_X1    g241(.A(new_n407_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n428_), .B1(new_n413_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n406_), .A2(KEYINPUT102), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT102), .B1(new_n406_), .B2(new_n445_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n442_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n450_), .A2(KEYINPUT103), .A3(new_n446_), .A4(new_n444_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n429_), .A2(KEYINPUT33), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n411_), .A2(new_n414_), .A3(new_n454_), .A4(new_n428_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT101), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(new_n328_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n322_), .A2(KEYINPUT101), .A3(new_n327_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n441_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n392_), .A2(new_n393_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT105), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n317_), .A2(new_n287_), .A3(new_n321_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n286_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n458_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n452_), .A2(new_n456_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n460_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n438_), .A2(new_n440_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n435_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n462_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT105), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n392_), .A2(new_n393_), .A3(new_n435_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n332_), .A2(new_n474_), .A3(new_n395_), .A4(new_n402_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n463_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n436_), .B1(new_n476_), .B2(new_n282_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G113gat), .B(G141gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT84), .ZN(new_n479_));
  XOR2_X1   g278(.A(G169gat), .B(G197gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G229gat), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G29gat), .B(G36gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G43gat), .B(G50gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n484_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G8gat), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n491_), .A2(KEYINPUT78), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493_));
  INV_X1    g292(.A(G1gat), .ZN(new_n494_));
  INV_X1    g293(.A(G8gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(KEYINPUT78), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n492_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n498_), .B1(new_n492_), .B2(new_n499_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n490_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n492_), .A2(new_n499_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n497_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n490_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n500_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n503_), .A2(KEYINPUT81), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT81), .B1(new_n503_), .B2(new_n507_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n483_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT82), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT82), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n513_), .B(new_n483_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n505_), .A2(new_n500_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(new_n490_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n490_), .B(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n518_), .B2(new_n515_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n482_), .B(KEYINPUT83), .Z(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n481_), .B1(new_n512_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT85), .ZN(new_n524_));
  INV_X1    g323(.A(new_n481_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n511_), .A2(new_n514_), .A3(new_n521_), .A4(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(KEYINPUT85), .B(new_n481_), .C1(new_n512_), .C2(new_n522_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT13), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G120gat), .B(G148gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT5), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G176gat), .B(G204gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G230gat), .A2(G233gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(G64gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(G57gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n421_), .A2(G64gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(KEYINPUT11), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT11), .B1(new_n539_), .B2(new_n540_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT67), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n543_), .A2(KEYINPUT67), .A3(new_n544_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n542_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n545_), .A3(new_n541_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G85gat), .B(G92gat), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT65), .ZN(new_n554_));
  AND3_X1   g353(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(KEYINPUT65), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT64), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n567_));
  NOR2_X1   g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n564_), .B(new_n565_), .C1(G99gat), .C2(G106gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n553_), .B1(new_n563_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT8), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT66), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n557_), .A2(new_n562_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n575_), .B(KEYINPUT8), .C1(new_n576_), .C2(new_n553_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n555_), .A2(new_n556_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(new_n573_), .A3(new_n552_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n574_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT10), .B(G99gat), .Z(new_n582_));
  INV_X1    g381(.A(G106gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n552_), .A2(KEYINPUT9), .ZN(new_n585_));
  INV_X1    g384(.A(G92gat), .ZN(new_n586_));
  OR3_X1    g385(.A1(new_n415_), .A2(new_n586_), .A3(KEYINPUT9), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n584_), .A2(new_n585_), .A3(new_n587_), .A4(new_n578_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n551_), .B1(new_n581_), .B2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n589_), .A2(KEYINPUT68), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n581_), .A2(new_n588_), .A3(new_n551_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n591_), .B1(new_n589_), .B2(KEYINPUT68), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n537_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n594_));
  INV_X1    g393(.A(new_n588_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n577_), .A2(new_n580_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n596_), .B2(new_n574_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n594_), .B1(new_n597_), .B2(new_n551_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n581_), .A2(new_n588_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n551_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(KEYINPUT12), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n598_), .A2(new_n536_), .A3(new_n591_), .A4(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n535_), .B1(new_n593_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n593_), .A2(new_n602_), .A3(new_n535_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n530_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n605_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n607_), .A2(KEYINPUT13), .A3(new_n603_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n609_), .A2(KEYINPUT69), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(KEYINPUT69), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n477_), .A2(new_n529_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n618_));
  AOI22_X1  g417(.A1(new_n597_), .A2(new_n506_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n599_), .A2(new_n518_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT73), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n617_), .A2(new_n618_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n619_), .B(new_n620_), .C1(new_n621_), .C2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n617_), .A2(new_n618_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n621_), .B(new_n625_), .C1(new_n599_), .C2(new_n490_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n599_), .B2(new_n490_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n518_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n597_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n626_), .B(new_n622_), .C1(new_n627_), .C2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT75), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n624_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT74), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(KEYINPUT36), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n624_), .A2(new_n630_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n636_), .A2(KEYINPUT36), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n637_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n624_), .A2(new_n630_), .A3(new_n631_), .A4(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n638_), .A2(new_n641_), .A3(KEYINPUT37), .A4(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT76), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n632_), .A2(new_n637_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT76), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(KEYINPUT37), .A4(new_n643_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n638_), .A2(new_n643_), .A3(new_n641_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT77), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n650_), .A2(KEYINPUT77), .A3(new_n651_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n649_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n515_), .B(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(new_n600_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n600_), .ZN(new_n660_));
  XOR2_X1   g459(.A(G127gat), .B(G155gat), .Z(new_n661_));
  XNOR2_X1  g460(.A(G183gat), .B(G211gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT17), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n659_), .A2(new_n660_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT79), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n665_), .A2(new_n669_), .A3(new_n666_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n668_), .B(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n656_), .A2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n613_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n494_), .A3(new_n435_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT38), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n650_), .B(KEYINPUT108), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n477_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n612_), .A2(new_n529_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n671_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G1gat), .B1(new_n681_), .B2(new_n437_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n675_), .A2(new_n682_), .ZN(G1324gat));
  AND2_X1   g482(.A1(new_n332_), .A2(new_n402_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n395_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n673_), .A2(new_n495_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n685_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G8gat), .B1(new_n681_), .B2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT39), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT39), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n692_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n686_), .B(new_n694_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1325gat));
  OAI21_X1  g495(.A(G15gat), .B1(new_n681_), .B2(new_n282_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(KEYINPUT41), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(KEYINPUT41), .ZN(new_n699_));
  INV_X1    g498(.A(new_n282_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n673_), .A2(new_n270_), .A3(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(new_n699_), .A3(new_n701_), .ZN(G1326gat));
  OAI21_X1  g501(.A(G22gat), .B1(new_n681_), .B2(new_n394_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT42), .ZN(new_n704_));
  INV_X1    g503(.A(G22gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n673_), .A2(new_n705_), .A3(new_n462_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1327gat));
  NOR2_X1   g506(.A1(new_n676_), .A2(new_n680_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n613_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G29gat), .B1(new_n710_), .B2(new_n435_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n649_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n477_), .A2(KEYINPUT43), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n475_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n715_));
  AOI211_X1 g514(.A(KEYINPUT105), .B(new_n462_), .C1(new_n468_), .C2(new_n470_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n282_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n436_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n714_), .B1(new_n719_), .B2(new_n656_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n679_), .B(new_n671_), .C1(new_n713_), .C2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n723_), .A2(G29gat), .A3(new_n435_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT43), .B1(new_n477_), .B2(new_n712_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n719_), .A2(new_n714_), .A3(new_n656_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n727_), .A2(KEYINPUT44), .A3(new_n679_), .A4(new_n671_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n711_), .B1(new_n724_), .B2(new_n728_), .ZN(G1328gat));
  NAND3_X1  g528(.A1(new_n723_), .A2(new_n685_), .A3(new_n728_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G36gat), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n613_), .A2(new_n732_), .A3(new_n685_), .A4(new_n708_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT45), .ZN(new_n734_));
  NOR2_X1   g533(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n731_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n687_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n732_), .B1(new_n738_), .B2(new_n728_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n733_), .B(KEYINPUT45), .Z(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1329gat));
  NAND4_X1  g541(.A1(new_n723_), .A2(G43gat), .A3(new_n700_), .A4(new_n728_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n267_), .B1(new_n709_), .B2(new_n282_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT47), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n743_), .A2(new_n747_), .A3(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1330gat));
  OR3_X1    g548(.A1(new_n709_), .A2(G50gat), .A3(new_n394_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n723_), .A2(new_n462_), .A3(new_n728_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT111), .ZN(new_n752_));
  OAI21_X1  g551(.A(G50gat), .B1(new_n751_), .B2(KEYINPUT111), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1331gat));
  AND2_X1   g553(.A1(new_n672_), .A2(new_n612_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n755_), .A2(KEYINPUT112), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n719_), .A3(new_n529_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(KEYINPUT112), .B2(new_n755_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n421_), .A3(new_n435_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n612_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n529_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n671_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n678_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G57gat), .B1(new_n764_), .B2(new_n437_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n759_), .A2(new_n765_), .ZN(G1332gat));
  AOI21_X1  g565(.A(new_n538_), .B1(new_n763_), .B2(new_n685_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT48), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n758_), .A2(new_n538_), .A3(new_n685_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1333gat));
  INV_X1    g569(.A(G71gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n763_), .B2(new_n700_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT49), .Z(new_n773_));
  NAND3_X1  g572(.A1(new_n758_), .A2(new_n771_), .A3(new_n700_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1334gat));
  INV_X1    g574(.A(G78gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n758_), .A2(new_n776_), .A3(new_n462_), .ZN(new_n777_));
  OAI21_X1  g576(.A(G78gat), .B1(new_n764_), .B2(new_n394_), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n778_), .A2(new_n779_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n777_), .A2(new_n780_), .A3(new_n781_), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n760_), .A2(new_n761_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n708_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n719_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n415_), .A3(new_n435_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n727_), .A2(new_n671_), .A3(new_n783_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G85gat), .B1(new_n788_), .B2(new_n437_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1336gat));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n586_), .A3(new_n685_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G92gat), .B1(new_n788_), .B2(new_n687_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n788_), .B2(new_n282_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n700_), .A2(new_n582_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n785_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g596(.A1(new_n786_), .A2(new_n583_), .A3(new_n462_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n727_), .A2(new_n462_), .A3(new_n671_), .A4(new_n783_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(new_n800_), .A3(G106gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n799_), .B2(G106gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT53), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n798_), .B(new_n805_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1339gat));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n508_), .A2(new_n509_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n520_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n519_), .A2(new_n810_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n481_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n526_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n815_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n816_), .A2(new_n817_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n591_), .B1(new_n589_), .B2(KEYINPUT12), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n594_), .B(new_n551_), .C1(new_n581_), .C2(new_n588_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n537_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n820_), .A2(new_n537_), .A3(new_n821_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(KEYINPUT55), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT115), .B1(new_n602_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(new_n827_), .A3(KEYINPUT55), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n824_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n819_), .B1(new_n829_), .B2(new_n535_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n826_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n602_), .A2(new_n825_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n832_), .A2(new_n822_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n534_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n607_), .B1(new_n830_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n818_), .B1(new_n836_), .B2(new_n761_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n808_), .B1(new_n837_), .B2(new_n677_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n529_), .B(new_n607_), .C1(new_n830_), .C2(new_n835_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT57), .B(new_n676_), .C1(new_n839_), .C2(new_n818_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n816_), .A2(new_n817_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n834_), .B2(new_n534_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n819_), .B(new_n535_), .C1(new_n831_), .C2(new_n833_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n605_), .B(new_n841_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n836_), .A2(KEYINPUT58), .A3(new_n841_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n656_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n838_), .A2(new_n840_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n671_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n671_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n851_), .B(KEYINPUT114), .C1(new_n606_), .C2(new_n608_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n712_), .A2(new_n852_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n712_), .A2(KEYINPUT54), .A3(new_n852_), .A4(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n850_), .A2(new_n861_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n282_), .A2(new_n403_), .A3(new_n437_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n761_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n862_), .A2(KEYINPUT59), .A3(new_n863_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT59), .B1(new_n862_), .B2(new_n863_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n529_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n867_), .B1(new_n872_), .B2(new_n866_), .ZN(G1340gat));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n874_));
  AOI21_X1  g673(.A(G120gat), .B1(new_n612_), .B2(new_n874_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n875_), .A2(KEYINPUT117), .B1(new_n874_), .B2(G120gat), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n865_), .B(new_n876_), .C1(KEYINPUT117), .C2(new_n875_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n760_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n878_));
  INV_X1    g677(.A(G120gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(G1341gat));
  AOI21_X1  g679(.A(G127gat), .B1(new_n865_), .B2(new_n680_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n869_), .A2(new_n871_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n680_), .A2(G127gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT118), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n881_), .B1(new_n882_), .B2(new_n884_), .ZN(G1342gat));
  OAI211_X1 g684(.A(G134gat), .B(new_n656_), .C1(new_n868_), .C2(new_n870_), .ZN(new_n886_));
  INV_X1    g685(.A(G134gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n864_), .B2(new_n676_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  OAI211_X1 g689(.A(KEYINPUT119), .B(new_n887_), .C1(new_n864_), .C2(new_n676_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n886_), .A2(new_n890_), .A3(new_n891_), .ZN(G1343gat));
  NOR4_X1   g691(.A1(new_n700_), .A2(new_n685_), .A3(new_n437_), .A4(new_n394_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n862_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n529_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT120), .B(G141gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1344gat));
  NOR2_X1   g696(.A1(new_n894_), .A2(new_n760_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n354_), .ZN(G1345gat));
  NOR2_X1   g698(.A1(new_n894_), .A2(new_n671_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT61), .B(G155gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903_));
  OAI21_X1  g702(.A(G162gat), .B1(new_n894_), .B2(new_n712_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n894_), .A2(G162gat), .A3(new_n676_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n903_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n906_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(KEYINPUT121), .A3(new_n904_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1347gat));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n860_), .B1(new_n849_), .B2(new_n671_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n700_), .A2(new_n685_), .A3(new_n437_), .A4(new_n394_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n761_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n911_), .B1(new_n915_), .B2(G169gat), .ZN(new_n916_));
  AOI211_X1 g715(.A(KEYINPUT62), .B(new_n227_), .C1(new_n914_), .C2(new_n761_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n913_), .ZN(new_n918_));
  AOI21_X1  g717(.A(KEYINPUT122), .B1(new_n862_), .B2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n912_), .A2(new_n920_), .A3(new_n913_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n761_), .A2(new_n311_), .ZN(new_n923_));
  OAI22_X1  g722(.A1(new_n916_), .A2(new_n917_), .B1(new_n922_), .B2(new_n923_), .ZN(G1348gat));
  NOR4_X1   g723(.A1(new_n912_), .A2(new_n222_), .A3(new_n760_), .A4(new_n913_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n862_), .A2(KEYINPUT122), .A3(new_n918_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n920_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n760_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT123), .B1(new_n928_), .B2(new_n226_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n612_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n930_), .A2(new_n931_), .A3(new_n310_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n925_), .B1(new_n929_), .B2(new_n932_), .ZN(G1349gat));
  AOI21_X1  g732(.A(G183gat), .B1(new_n914_), .B2(new_n680_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n671_), .A2(new_n258_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(KEYINPUT124), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n938_), .B(new_n935_), .C1(new_n919_), .C2(new_n921_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n934_), .B1(new_n937_), .B2(new_n939_), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n922_), .B2(new_n712_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n677_), .A2(new_n259_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n922_), .B2(new_n942_), .ZN(G1351gat));
  NAND3_X1  g742(.A1(new_n282_), .A2(new_n437_), .A3(new_n462_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n685_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n945_), .B2(new_n944_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n862_), .A2(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n529_), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT126), .B(G197gat), .Z(new_n950_));
  XNOR2_X1  g749(.A(new_n949_), .B(new_n950_), .ZN(G1352gat));
  INV_X1    g750(.A(new_n948_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n612_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n948_), .A2(new_n671_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n955_), .B1(new_n956_), .B2(new_n958_), .ZN(new_n959_));
  OAI211_X1 g758(.A(KEYINPUT127), .B(new_n957_), .C1(new_n948_), .C2(new_n671_), .ZN(new_n960_));
  XOR2_X1   g759(.A(KEYINPUT63), .B(G211gat), .Z(new_n961_));
  AOI22_X1  g760(.A1(new_n959_), .A2(new_n960_), .B1(new_n956_), .B2(new_n961_), .ZN(G1354gat));
  OR3_X1    g761(.A1(new_n948_), .A2(G218gat), .A3(new_n676_), .ZN(new_n963_));
  OAI21_X1  g762(.A(G218gat), .B1(new_n948_), .B2(new_n712_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1355gat));
endmodule


