//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n978_, new_n979_, new_n980_, new_n982_, new_n983_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n990_, new_n991_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n998_, new_n999_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(G230gat), .ZN(new_n203_));
  INV_X1    g002(.A(G233gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207_));
  INV_X1    g006(.A(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT7), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n217_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n211_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G85gat), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(KEYINPUT8), .A3(new_n224_), .ZN(new_n228_));
  OR2_X1    g027(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n229_), .A2(KEYINPUT64), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT64), .B1(new_n229_), .B2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n209_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n222_), .A2(KEYINPUT9), .A3(new_n223_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n223_), .A2(KEYINPUT9), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n216_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n227_), .A2(new_n228_), .A3(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G64gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G78gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(KEYINPUT11), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n242_));
  INV_X1    g041(.A(new_n240_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n241_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n238_), .A2(new_n247_), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n225_), .A2(new_n226_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n228_), .A3(new_n246_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n206_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AOI211_X1 g052(.A(KEYINPUT66), .B(new_n206_), .C1(new_n248_), .C2(new_n250_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n206_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT12), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n246_), .B1(new_n249_), .B2(new_n228_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(KEYINPUT67), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n248_), .A2(new_n260_), .A3(KEYINPUT12), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n256_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G120gat), .B(G148gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n255_), .A2(new_n262_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  AND4_X1   g068(.A1(new_n228_), .A2(new_n227_), .A3(new_n237_), .A4(new_n246_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n205_), .B1(new_n258_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT66), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n251_), .A2(new_n252_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n256_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT12), .B1(new_n248_), .B2(new_n260_), .ZN(new_n276_));
  AOI211_X1 g075(.A(KEYINPUT67), .B(new_n257_), .C1(new_n238_), .C2(new_n247_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n269_), .B1(new_n274_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n202_), .B1(new_n268_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n267_), .B1(new_n255_), .B2(new_n262_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n274_), .A2(new_n278_), .A3(new_n269_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(KEYINPUT13), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT69), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n291_));
  NAND2_X1  g090(.A1(G232gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G43gat), .B(G50gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G36gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G29gat), .ZN(new_n297_));
  INV_X1    g096(.A(G29gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G36gat), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n297_), .A2(new_n299_), .A3(KEYINPUT71), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT71), .B1(new_n297_), .B2(new_n299_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n295_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n299_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n297_), .A2(new_n299_), .A3(KEYINPUT71), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(new_n294_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n302_), .A2(new_n307_), .A3(KEYINPUT15), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n228_), .A2(new_n249_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n238_), .A2(new_n308_), .ZN(new_n313_));
  OAI211_X1 g112(.A(KEYINPUT35), .B(new_n293_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G190gat), .B(G218gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G134gat), .B(G162gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(KEYINPUT36), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n310_), .A2(new_n311_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n238_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n293_), .A2(KEYINPUT35), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n293_), .A2(KEYINPUT35), .ZN(new_n322_));
  INV_X1    g121(.A(new_n308_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n249_), .A2(new_n323_), .A3(new_n228_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n314_), .A2(new_n318_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT72), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n314_), .A2(new_n328_), .A3(new_n325_), .A4(new_n318_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT37), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n314_), .A2(new_n325_), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n317_), .B(KEYINPUT36), .Z(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n333_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n330_), .B(new_n331_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n334_), .B(KEYINPUT73), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n330_), .A2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n337_), .B(KEYINPUT75), .C1(new_n340_), .C2(new_n331_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n336_), .A2(new_n335_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(new_n331_), .A4(new_n330_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT14), .ZN(new_n348_));
  INV_X1    g147(.A(G8gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT76), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G8gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n348_), .B1(new_n353_), .B2(G1gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(G15gat), .B(G22gat), .Z(new_n355_));
  OAI21_X1  g154(.A(new_n347_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT76), .B(G8gat), .ZN(new_n357_));
  INV_X1    g156(.A(G1gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT14), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n355_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(KEYINPUT77), .A3(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G1gat), .B(G8gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n356_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n356_), .B2(new_n361_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G127gat), .B(G155gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT16), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G183gat), .B(G211gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT16), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n368_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT17), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G231gat), .A2(G233gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(KEYINPUT78), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n377_), .B2(KEYINPUT78), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n246_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n377_), .A2(KEYINPUT78), .ZN(new_n383_));
  INV_X1    g182(.A(new_n378_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n247_), .B1(new_n385_), .B2(new_n379_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n367_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n246_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n379_), .A3(new_n247_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n366_), .A3(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n376_), .A2(KEYINPUT17), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n387_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n346_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n290_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n396_), .B(G15gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT30), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G71gat), .B(G99gat), .ZN(new_n399_));
  INV_X1    g198(.A(G43gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OR3_X1    g201(.A1(KEYINPUT85), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT85), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(G169gat), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n404_), .ZN(new_n406_));
  INV_X1    g205(.A(G169gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G183gat), .ZN(new_n409_));
  INV_X1    g208(.A(G190gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT23), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT23), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(G183gat), .A3(G190gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n415_));
  OR2_X1    g214(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n410_), .A3(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n414_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n414_), .B2(new_n418_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n405_), .B(new_n408_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT24), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT24), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(new_n426_), .B2(new_n422_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n411_), .A2(KEYINPUT84), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n429_), .B(KEYINPUT23), .C1(new_n409_), .C2(new_n410_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n431_), .B2(new_n413_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G190gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT26), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n437_));
  NOR2_X1   g236(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n438_));
  OAI21_X1  g237(.A(G183gat), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(KEYINPUT82), .B(G183gat), .C1(new_n437_), .C2(new_n438_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n416_), .A2(KEYINPUT25), .A3(new_n417_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n436_), .A2(new_n441_), .A3(new_n442_), .A4(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n432_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n402_), .B1(new_n421_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n421_), .A2(new_n445_), .A3(new_n402_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n398_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n398_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n446_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT88), .B1(new_n449_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G127gat), .B(G134gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G113gat), .B(G120gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT31), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n447_), .A2(new_n398_), .A3(new_n448_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n451_), .B1(new_n450_), .B2(new_n446_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT87), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n453_), .B(new_n457_), .C1(new_n460_), .C2(KEYINPUT88), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n462_));
  INV_X1    g261(.A(new_n457_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n449_), .A2(new_n452_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n462_), .B(new_n463_), .C1(new_n464_), .C2(KEYINPUT87), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT99), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n407_), .A2(KEYINPUT22), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT22), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G169gat), .ZN(new_n471_));
  INV_X1    g270(.A(G176gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT95), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n425_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n473_), .B2(new_n425_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n413_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(G183gat), .A2(G190gat), .ZN(new_n479_));
  OAI22_X1  g278(.A1(new_n475_), .A2(new_n476_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n427_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT25), .B(G183gat), .Z(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT26), .B(G190gat), .Z(new_n483_));
  OAI211_X1 g282(.A(new_n481_), .B(new_n414_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(G197gat), .A2(G204gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G197gat), .A2(G204gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT21), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(KEYINPUT21), .A3(new_n487_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G211gat), .B(G218gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n491_), .A2(new_n492_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n468_), .B1(new_n485_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G226gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT19), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n493_), .A2(new_n494_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n421_), .A2(new_n445_), .A3(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n496_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n480_), .A2(new_n500_), .A3(new_n484_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT20), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT98), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n500_), .B1(new_n421_), .B2(new_n445_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT98), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n508_), .A3(KEYINPUT20), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n502_), .B1(new_n510_), .B2(new_n498_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G8gat), .B(G36gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n467_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n485_), .A2(new_n495_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(KEYINPUT20), .A3(new_n501_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n498_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n507_), .A2(KEYINPUT20), .A3(new_n499_), .A4(new_n503_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT27), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n516_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n506_), .B1(new_n504_), .B2(KEYINPUT98), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n499_), .B1(new_n526_), .B2(new_n509_), .ZN(new_n527_));
  OAI211_X1 g326(.A(KEYINPUT99), .B(new_n525_), .C1(new_n527_), .C2(new_n502_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n517_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G225gat), .A2(G233gat), .ZN(new_n530_));
  INV_X1    g329(.A(G155gat), .ZN(new_n531_));
  INV_X1    g330(.A(G162gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT89), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(G155gat), .B2(G162gat), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n533_), .B(new_n535_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n537_), .A2(KEYINPUT90), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(KEYINPUT90), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT3), .ZN(new_n541_));
  INV_X1    g340(.A(G141gat), .ZN(new_n542_));
  INV_X1    g341(.A(G148gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G141gat), .A2(G148gat), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT2), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n536_), .B1(new_n540_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT1), .B1(new_n531_), .B2(new_n532_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT1), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(G155gat), .A3(G162gat), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n552_), .A2(new_n533_), .A3(new_n535_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n542_), .A2(new_n543_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n545_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n456_), .B1(new_n551_), .B2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n454_), .B(new_n455_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(new_n556_), .A3(new_n545_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n549_), .B1(new_n539_), .B2(new_n538_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n559_), .B(new_n560_), .C1(new_n561_), .C2(new_n536_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(KEYINPUT4), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT4), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n564_), .B(new_n456_), .C1(new_n551_), .C2(new_n557_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n530_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G1gat), .B(G29gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G85gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT0), .B(G57gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n530_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n566_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n571_), .B1(new_n566_), .B2(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT91), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n551_), .A2(new_n557_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT29), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT28), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT28), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n579_), .A2(new_n583_), .A3(new_n580_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G22gat), .B(G50gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n585_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n578_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(KEYINPUT91), .A3(new_n586_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n495_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n592_));
  OR2_X1    g391(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(G233gat), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n495_), .B2(KEYINPUT93), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  OAI221_X1 g396(.A(new_n495_), .B1(KEYINPUT93), .B2(new_n595_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G78gat), .B(G106gat), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n600_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n589_), .A2(new_n591_), .A3(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n587_), .A2(new_n588_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(KEYINPUT94), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n597_), .A2(new_n598_), .A3(new_n608_), .A4(new_n602_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n606_), .A2(new_n607_), .A3(new_n601_), .A4(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n577_), .B1(new_n605_), .B2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n499_), .B1(new_n496_), .B2(new_n501_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n504_), .A2(new_n506_), .A3(new_n498_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n525_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT27), .B1(new_n614_), .B2(new_n522_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n529_), .A2(new_n611_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n558_), .A2(new_n572_), .A3(new_n562_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(new_n570_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n563_), .A2(new_n530_), .A3(new_n565_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n618_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n620_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n614_), .B(new_n522_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n576_), .A2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT33), .B(new_n571_), .C1(new_n566_), .C2(new_n573_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n516_), .A2(KEYINPUT32), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n510_), .A2(new_n498_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n502_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n520_), .A2(new_n521_), .A3(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n563_), .A2(new_n565_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n572_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n573_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n570_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n633_), .B1(new_n637_), .B2(new_n574_), .ZN(new_n638_));
  OAI22_X1  g437(.A1(new_n624_), .A2(new_n628_), .B1(new_n632_), .B2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n605_), .A2(new_n610_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n466_), .B1(new_n617_), .B2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n637_), .A2(new_n574_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n461_), .A2(new_n643_), .A3(new_n465_), .ZN(new_n644_));
  AND4_X1   g443(.A1(new_n640_), .A2(new_n644_), .A3(new_n616_), .A4(new_n529_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n647_), .B(new_n648_), .Z(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(KEYINPUT79), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n356_), .A2(new_n361_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n362_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n319_), .A2(new_n363_), .A3(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n323_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(G229gat), .A2(G233gat), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(new_n308_), .A3(new_n363_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n650_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n656_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n364_), .A2(new_n365_), .A3(new_n323_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n308_), .B1(new_n653_), .B2(new_n363_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n664_), .B(new_n665_), .C1(KEYINPUT79), .C2(new_n649_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n660_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n646_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n395_), .A2(new_n669_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n670_), .A2(G1gat), .A3(new_n643_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(KEYINPUT38), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT102), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n342_), .A2(new_n330_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n646_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n393_), .A2(new_n667_), .A3(new_n280_), .A4(new_n283_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT101), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G1gat), .B1(new_n679_), .B2(new_n643_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n671_), .A2(KEYINPUT38), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(KEYINPUT100), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n681_), .A2(KEYINPUT100), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n673_), .B(new_n680_), .C1(new_n682_), .C2(new_n683_), .ZN(G1324gat));
  OAI21_X1  g483(.A(new_n525_), .B1(new_n527_), .B2(new_n502_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n523_), .B1(new_n685_), .B2(new_n467_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n615_), .B1(new_n686_), .B2(new_n528_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G8gat), .B1(new_n679_), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT39), .ZN(new_n689_));
  INV_X1    g488(.A(new_n687_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n357_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n670_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1325gat));
  INV_X1    g493(.A(new_n466_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G15gat), .B1(new_n679_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT41), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n670_), .A2(G15gat), .A3(new_n695_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1326gat));
  OAI21_X1  g498(.A(G22gat), .B1(new_n679_), .B2(new_n640_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT42), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n640_), .A2(G22gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n670_), .B2(new_n702_), .ZN(G1327gat));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n646_), .B2(new_n346_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n706_), .B(new_n345_), .C1(new_n642_), .C2(new_n645_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n284_), .A2(new_n668_), .A3(new_n393_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n704_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n708_), .A2(KEYINPUT104), .A3(KEYINPUT44), .A4(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n710_), .A2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n643_), .A2(new_n298_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n714_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n675_), .A2(new_n392_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(new_n284_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n669_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G29gat), .B1(new_n722_), .B2(new_n577_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n718_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT105), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n718_), .A2(new_n727_), .A3(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(KEYINPUT46), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n716_), .A2(new_n690_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n296_), .B1(new_n733_), .B2(new_n714_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n690_), .A2(new_n296_), .ZN(new_n735_));
  OR3_X1    g534(.A1(new_n721_), .A2(KEYINPUT106), .A3(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT106), .B1(new_n721_), .B2(new_n735_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n736_), .A2(KEYINPUT45), .A3(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n731_), .B1(new_n734_), .B2(new_n742_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n736_), .A2(KEYINPUT45), .A3(new_n737_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT45), .B1(new_n736_), .B2(new_n737_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n731_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n732_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n746_), .B(new_n747_), .C1(new_n748_), .C2(new_n296_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n743_), .A2(new_n749_), .ZN(G1329gat));
  NOR2_X1   g549(.A1(new_n695_), .A2(new_n400_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n714_), .A2(new_n716_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G43gat), .B1(new_n722_), .B2(new_n466_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(new_n754_), .A3(new_n756_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1330gat));
  OR3_X1    g559(.A1(new_n721_), .A2(G50gat), .A3(new_n640_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n640_), .B1(new_n710_), .B2(new_n715_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n714_), .A2(KEYINPUT109), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G50gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT109), .B1(new_n714_), .B2(new_n762_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(G1331gat));
  NOR2_X1   g565(.A1(new_n392_), .A2(new_n667_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n676_), .A2(new_n290_), .A3(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(G57gat), .A3(new_n577_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT111), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT110), .B1(new_n646_), .B2(new_n667_), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n687_), .A2(new_n611_), .B1(new_n640_), .B2(new_n639_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n687_), .A2(new_n640_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n644_), .ZN(new_n774_));
  OAI22_X1  g573(.A1(new_n772_), .A2(new_n466_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n668_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n771_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n394_), .A2(new_n285_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G57gat), .B1(new_n781_), .B2(new_n577_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n770_), .A2(new_n782_), .ZN(G1332gat));
  OR3_X1    g582(.A1(new_n780_), .A2(G64gat), .A3(new_n687_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n768_), .A2(new_n690_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(G64gat), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(KEYINPUT48), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(KEYINPUT48), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(G1333gat));
  OR3_X1    g588(.A1(new_n780_), .A2(G71gat), .A3(new_n695_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n768_), .A2(new_n466_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G71gat), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(KEYINPUT49), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(KEYINPUT49), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(G1334gat));
  OR3_X1    g594(.A1(new_n780_), .A2(G78gat), .A3(new_n640_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n640_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n768_), .A2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(G78gat), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G78gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n796_), .B1(new_n800_), .B2(new_n801_), .ZN(G1335gat));
  NOR2_X1   g601(.A1(new_n289_), .A2(new_n719_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n778_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT113), .B1(new_n778_), .B2(new_n803_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(new_n220_), .A3(new_n577_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n285_), .A2(new_n667_), .A3(new_n393_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n708_), .A2(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(new_n577_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n810_), .B1(new_n220_), .B2(new_n813_), .ZN(G1336gat));
  NAND3_X1  g613(.A1(new_n809_), .A2(new_n221_), .A3(new_n690_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n812_), .A2(new_n690_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n221_), .B2(new_n816_), .ZN(G1337gat));
  OAI21_X1  g616(.A(new_n466_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n812_), .A2(new_n466_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n808_), .A2(new_n818_), .B1(new_n208_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g620(.A(new_n209_), .B(new_n797_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n706_), .B1(new_n775_), .B2(new_n345_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n707_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n797_), .B(new_n811_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n708_), .A2(KEYINPUT114), .A3(new_n797_), .A4(new_n811_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n209_), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n823_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n823_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n831_), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n833_), .B(new_n834_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n822_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT53), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n822_), .B(new_n838_), .C1(new_n832_), .C2(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1339gat));
  INV_X1    g639(.A(G113gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n668_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n656_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n654_), .A2(new_n655_), .A3(new_n661_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n649_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n649_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT118), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n844_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n661_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n846_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n649_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n851_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n848_), .A2(new_n854_), .A3(new_n282_), .ZN(new_n855_));
  AND2_X1   g654(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT55), .B(new_n275_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n278_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n250_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n205_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n259_), .A2(new_n261_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n864_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n275_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n859_), .A2(new_n861_), .A3(new_n863_), .A4(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n267_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n856_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n866_), .B(new_n267_), .C1(KEYINPUT119), .C2(KEYINPUT56), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n855_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n345_), .B1(new_n871_), .B2(KEYINPUT58), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873_));
  AOI211_X1 g672(.A(new_n873_), .B(new_n855_), .C1(new_n869_), .C2(new_n870_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n268_), .A2(new_n279_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n848_), .A2(new_n854_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n667_), .A2(new_n282_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT56), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT117), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n867_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n882_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n866_), .A2(new_n267_), .A3(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n879_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n876_), .B1(new_n886_), .B2(new_n675_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n866_), .A2(new_n267_), .A3(new_n884_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n884_), .B1(new_n866_), .B2(new_n267_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n880_), .ZN(new_n890_));
  OAI211_X1 g689(.A(KEYINPUT57), .B(new_n674_), .C1(new_n890_), .C2(new_n879_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n887_), .A2(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n392_), .B1(new_n875_), .B2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n767_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT54), .B1(new_n345_), .B2(new_n894_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n767_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n341_), .A4(new_n344_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n895_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n893_), .A2(new_n900_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n773_), .A2(new_n695_), .A3(new_n643_), .ZN(new_n902_));
  AOI21_X1  g701(.A(KEYINPUT59), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n887_), .B(new_n891_), .C1(new_n872_), .C2(new_n874_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n899_), .B1(new_n904_), .B2(new_n392_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906_));
  INV_X1    g705(.A(new_n902_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n842_), .B1(new_n903_), .B2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n893_), .B2(new_n900_), .ZN(new_n910_));
  AOI211_X1 g709(.A(KEYINPUT120), .B(G113gat), .C1(new_n910_), .C2(new_n667_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n887_), .A2(new_n891_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n869_), .A2(new_n870_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n873_), .B1(new_n914_), .B2(new_n855_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n871_), .A2(KEYINPUT58), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n345_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n393_), .B1(new_n913_), .B2(new_n917_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n667_), .B(new_n902_), .C1(new_n918_), .C2(new_n899_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n912_), .B1(new_n919_), .B2(new_n841_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n909_), .B1(new_n911_), .B2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT121), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n909_), .B(new_n923_), .C1(new_n911_), .C2(new_n920_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1340gat));
  INV_X1    g724(.A(G120gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n901_), .A2(KEYINPUT59), .A3(new_n902_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n906_), .B1(new_n905_), .B2(new_n907_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n926_), .B1(new_n929_), .B2(new_n290_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n910_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n926_), .B1(new_n285_), .B2(KEYINPUT60), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n932_), .B1(KEYINPUT60), .B2(new_n926_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT122), .B1(new_n930_), .B2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n289_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n937_));
  OAI221_X1 g736(.A(new_n936_), .B1(new_n931_), .B2(new_n933_), .C1(new_n937_), .C2(new_n926_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n935_), .A2(new_n938_), .ZN(G1341gat));
  NAND2_X1  g738(.A1(new_n393_), .A2(G127gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT123), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n941_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943_));
  AOI21_X1  g742(.A(G127gat), .B1(new_n910_), .B2(new_n393_), .ZN(new_n944_));
  OR3_X1    g743(.A1(new_n942_), .A2(new_n943_), .A3(new_n944_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n942_), .B2(new_n944_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1342gat));
  AOI21_X1  g746(.A(G134gat), .B1(new_n910_), .B2(new_n675_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n345_), .A2(G134gat), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(KEYINPUT125), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n948_), .B1(new_n929_), .B2(new_n950_), .ZN(G1343gat));
  NOR4_X1   g750(.A1(new_n690_), .A2(new_n640_), .A3(new_n466_), .A4(new_n643_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n901_), .A2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n953_), .A2(new_n668_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(new_n542_), .ZN(G1344gat));
  NOR2_X1   g754(.A1(new_n953_), .A2(new_n289_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(new_n543_), .ZN(G1345gat));
  NOR2_X1   g756(.A1(new_n953_), .A2(new_n392_), .ZN(new_n958_));
  XOR2_X1   g757(.A(KEYINPUT61), .B(G155gat), .Z(new_n959_));
  XNOR2_X1  g758(.A(new_n958_), .B(new_n959_), .ZN(G1346gat));
  OAI21_X1  g759(.A(new_n532_), .B1(new_n953_), .B2(new_n674_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(KEYINPUT126), .ZN(new_n962_));
  NOR3_X1   g761(.A1(new_n953_), .A2(new_n532_), .A3(new_n346_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1347gat));
  NOR2_X1   g763(.A1(new_n905_), .A2(new_n687_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n774_), .A2(new_n797_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G169gat), .B1(new_n967_), .B2(new_n668_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n967_), .ZN(new_n971_));
  NAND4_X1  g770(.A1(new_n971_), .A2(new_n667_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n972_));
  OAI211_X1 g771(.A(KEYINPUT62), .B(G169gat), .C1(new_n967_), .C2(new_n668_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n970_), .A2(new_n972_), .A3(new_n973_), .ZN(G1348gat));
  OAI21_X1  g773(.A(G176gat), .B1(new_n967_), .B2(new_n289_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n284_), .A2(new_n472_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n975_), .B1(new_n967_), .B2(new_n976_), .ZN(G1349gat));
  NOR2_X1   g776(.A1(new_n967_), .A2(new_n392_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n416_), .A2(new_n417_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n978_), .A2(new_n979_), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n980_), .B1(new_n482_), .B2(new_n978_), .ZN(G1350gat));
  OAI21_X1  g780(.A(G190gat), .B1(new_n967_), .B2(new_n346_), .ZN(new_n982_));
  OR2_X1    g781(.A1(new_n674_), .A2(new_n483_), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n982_), .B1(new_n967_), .B2(new_n983_), .ZN(G1351gat));
  NOR3_X1   g783(.A1(new_n466_), .A2(new_n640_), .A3(new_n577_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n965_), .A2(new_n985_), .ZN(new_n986_));
  INV_X1    g785(.A(new_n986_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n987_), .A2(new_n667_), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g788(.A1(new_n986_), .A2(new_n289_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(KEYINPUT127), .B(G204gat), .ZN(new_n991_));
  XNOR2_X1  g790(.A(new_n990_), .B(new_n991_), .ZN(G1353gat));
  NAND3_X1  g791(.A1(new_n965_), .A2(new_n393_), .A3(new_n985_), .ZN(new_n993_));
  NOR2_X1   g792(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n994_));
  AND2_X1   g793(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n995_));
  NOR3_X1   g794(.A1(new_n993_), .A2(new_n994_), .A3(new_n995_), .ZN(new_n996_));
  AOI21_X1  g795(.A(new_n996_), .B1(new_n993_), .B2(new_n994_), .ZN(G1354gat));
  OR3_X1    g796(.A1(new_n986_), .A2(G218gat), .A3(new_n674_), .ZN(new_n998_));
  OAI21_X1  g797(.A(G218gat), .B1(new_n986_), .B2(new_n346_), .ZN(new_n999_));
  NAND2_X1  g798(.A1(new_n998_), .A2(new_n999_), .ZN(G1355gat));
endmodule


