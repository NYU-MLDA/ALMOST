//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G29gat), .B(G36gat), .Z(new_n206_));
  XOR2_X1   g005(.A(G43gat), .B(G50gat), .Z(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  XOR2_X1   g007(.A(G1gat), .B(G8gat), .Z(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT75), .B(G15gat), .ZN(new_n211_));
  INV_X1    g010(.A(G22gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G1gat), .A2(G8gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT14), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n213_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(new_n213_), .B2(new_n216_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n210_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n219_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n209_), .A3(new_n217_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n208_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n208_), .B(KEYINPUT15), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n222_), .A3(new_n208_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n228_), .B1(new_n224_), .B2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n205_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n224_), .A2(new_n231_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n229_), .B(new_n204_), .C1(new_n234_), .C2(new_n228_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n235_), .A3(KEYINPUT82), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n237_), .B(new_n205_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G120gat), .B(G148gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT72), .ZN(new_n241_));
  XOR2_X1   g040(.A(G176gat), .B(G204gat), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT12), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT10), .B(G99gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT64), .ZN(new_n249_));
  INV_X1    g048(.A(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT65), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT6), .ZN(new_n255_));
  AND2_X1   g054(.A1(G99gat), .A2(G106gat), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n253_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G85gat), .A2(G92gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT9), .ZN(new_n261_));
  XOR2_X1   g060(.A(G85gat), .B(G92gat), .Z(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(KEYINPUT9), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n251_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n258_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n253_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT66), .B1(new_n257_), .B2(new_n258_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G99gat), .A2(G106gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT7), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n269_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n262_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT67), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(new_n276_), .A3(new_n262_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(KEYINPUT8), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n259_), .A2(new_n272_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT8), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n262_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n265_), .B1(new_n278_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G57gat), .B(G64gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n284_));
  XOR2_X1   g083(.A(G71gat), .B(G78gat), .Z(new_n285_));
  OR2_X1    g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n285_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n247_), .B1(new_n282_), .B2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(KEYINPUT69), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(KEYINPUT69), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT12), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n277_), .A2(KEYINPUT8), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n276_), .B1(new_n273_), .B2(new_n262_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n281_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n296_), .B2(new_n264_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G230gat), .A2(G233gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n282_), .A2(new_n289_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n290_), .A2(new_n298_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT70), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n296_), .A2(new_n264_), .A3(new_n289_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(new_n297_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n299_), .A4(new_n290_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n299_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n289_), .B1(new_n296_), .B2(new_n264_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(new_n303_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT68), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n246_), .B1(new_n307_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n310_), .B(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n314_), .A2(new_n302_), .A3(new_n306_), .A4(new_n245_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(KEYINPUT13), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT13), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n239_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT85), .ZN(new_n321_));
  INV_X1    g120(.A(G134gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G127gat), .ZN(new_n323_));
  INV_X1    g122(.A(G127gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G134gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G120gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G113gat), .ZN(new_n328_));
  INV_X1    g127(.A(G113gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G120gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n321_), .B1(new_n326_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n331_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n323_), .A2(new_n325_), .A3(new_n328_), .A4(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n335_), .B2(new_n321_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT31), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n337_), .A2(KEYINPUT86), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n337_), .A2(KEYINPUT86), .ZN(new_n339_));
  INV_X1    g138(.A(G183gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT25), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G183gat), .ZN(new_n343_));
  INV_X1    g142(.A(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT26), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G190gat), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n341_), .A2(new_n343_), .A3(new_n345_), .A4(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  OR3_X1    g151(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n353_));
  INV_X1    g152(.A(G169gat), .ZN(new_n354_));
  INV_X1    g153(.A(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(KEYINPUT24), .A3(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n348_), .A2(new_n352_), .A3(new_n353_), .A4(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G169gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n351_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n340_), .A2(new_n344_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(new_n349_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n359_), .A2(new_n365_), .A3(KEYINPUT83), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT83), .B1(new_n359_), .B2(new_n365_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT30), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT84), .B(G43gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(G15gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G71gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G99gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n371_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n371_), .A2(new_n378_), .ZN(new_n380_));
  AOI211_X1 g179(.A(new_n338_), .B(new_n339_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n379_), .A2(new_n338_), .A3(new_n380_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386_));
  OR2_X1    g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388_));
  INV_X1    g187(.A(G141gat), .ZN(new_n389_));
  INV_X1    g188(.A(G148gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT87), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(KEYINPUT87), .A3(new_n388_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n386_), .B(new_n387_), .C1(new_n396_), .C2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n386_), .A2(KEYINPUT1), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT1), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(G155gat), .A3(G162gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n406_), .A3(new_n387_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n394_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n397_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n385_), .B1(new_n403_), .B2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(G197gat), .A2(G204gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G197gat), .A2(G204gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT21), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(KEYINPUT21), .A3(new_n412_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G211gat), .B(G218gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n416_), .A2(new_n417_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(G228gat), .B(G233gat), .C1(new_n410_), .C2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n387_), .A2(new_n386_), .ZN(new_n423_));
  NOR4_X1   g222(.A1(new_n392_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT87), .B1(new_n394_), .B2(new_n388_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n402_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n409_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n422_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n403_), .A2(KEYINPUT88), .A3(new_n409_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(KEYINPUT29), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT90), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G228gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT89), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n420_), .A2(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n432_), .A2(new_n433_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n433_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n421_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n430_), .A2(new_n431_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT28), .B1(new_n440_), .B2(KEYINPUT29), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n430_), .A2(new_n431_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT28), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n385_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n439_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n444_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n446_), .B(new_n421_), .C1(new_n438_), .C2(new_n437_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G78gat), .B(G106gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(G22gat), .B(G50gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n445_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n402_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n409_), .B(new_n335_), .C1(new_n455_), .C2(new_n423_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT94), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT94), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n403_), .A2(new_n458_), .A3(new_n409_), .A4(new_n335_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n430_), .A2(new_n431_), .A3(new_n336_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G225gat), .A2(G233gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT96), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n460_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(G85gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT0), .B(G57gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n467_), .B(new_n468_), .Z(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n460_), .A2(KEYINPUT4), .A3(new_n461_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT95), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT95), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n460_), .A2(new_n461_), .A3(new_n473_), .A4(KEYINPUT4), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT4), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n440_), .A2(KEYINPUT97), .A3(new_n476_), .A4(new_n336_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT97), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n461_), .B2(KEYINPUT4), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n464_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n470_), .B1(new_n475_), .B2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n481_), .A2(KEYINPUT33), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G226gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT19), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n484_), .B(KEYINPUT91), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n359_), .A2(new_n365_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n359_), .A2(new_n365_), .A3(KEYINPUT83), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n420_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT20), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n418_), .A2(new_n419_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n486_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n491_), .B1(new_n490_), .B2(KEYINPUT20), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n485_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G8gat), .B(G36gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT18), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G64gat), .B(G92gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  OAI21_X1  g300(.A(new_n493_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n486_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n484_), .B1(new_n503_), .B2(new_n420_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n504_), .A3(KEYINPUT20), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n502_), .A2(new_n504_), .A3(KEYINPUT93), .A4(KEYINPUT20), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n497_), .A2(new_n501_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n501_), .B1(new_n497_), .B2(new_n509_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n475_), .A2(new_n480_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n465_), .A2(KEYINPUT33), .A3(new_n469_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n463_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n475_), .A2(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n460_), .A2(new_n461_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n469_), .B1(new_n517_), .B2(new_n463_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n513_), .A2(new_n514_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n482_), .A2(new_n512_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT101), .ZN(new_n521_));
  INV_X1    g320(.A(new_n470_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n513_), .B2(new_n522_), .ZN(new_n523_));
  AOI211_X1 g322(.A(KEYINPUT101), .B(new_n470_), .C1(new_n475_), .C2(new_n480_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n465_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n475_), .B2(new_n480_), .ZN(new_n526_));
  OAI22_X1  g325(.A1(new_n523_), .A2(new_n524_), .B1(new_n526_), .B2(new_n469_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n497_), .A2(new_n509_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n501_), .A2(KEYINPUT32), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n366_), .A2(new_n367_), .A3(new_n493_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT92), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n485_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n494_), .A4(new_n492_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT100), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n493_), .B1(KEYINPUT99), .B2(new_n486_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(KEYINPUT99), .B2(new_n486_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(KEYINPUT20), .A3(new_n502_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n535_), .A2(new_n536_), .B1(new_n484_), .B2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n495_), .A2(new_n496_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(KEYINPUT100), .A3(new_n534_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n530_), .B1(new_n529_), .B2(new_n543_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n520_), .A2(KEYINPUT98), .B1(new_n527_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT98), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n482_), .A2(new_n512_), .A3(new_n519_), .A4(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n454_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n501_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n501_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT27), .B1(new_n528_), .B2(new_n550_), .ZN(new_n551_));
  OAI22_X1  g350(.A1(new_n512_), .A2(KEYINPUT27), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n552_), .A2(new_n527_), .A3(new_n453_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n384_), .B1(new_n548_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n527_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n383_), .A2(new_n555_), .A3(new_n556_), .A4(new_n453_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n320_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT80), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n291_), .A2(new_n292_), .ZN(new_n561_));
  INV_X1    g360(.A(G231gat), .ZN(new_n562_));
  INV_X1    g361(.A(G233gat), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n220_), .A2(new_n222_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n561_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n220_), .A2(new_n222_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n561_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n220_), .A2(new_n222_), .A3(new_n564_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n567_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G127gat), .B(G155gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT79), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT79), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n574_), .A2(new_n584_), .A3(new_n581_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n289_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n289_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n570_), .A2(new_n588_), .A3(new_n572_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n579_), .B(KEYINPUT17), .Z(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n560_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  AOI211_X1 g392(.A(KEYINPUT80), .B(new_n593_), .C1(new_n583_), .C2(new_n585_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n559_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n585_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n584_), .B1(new_n574_), .B2(new_n581_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n591_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT80), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n586_), .A2(new_n560_), .A3(new_n591_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(KEYINPUT81), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT36), .Z(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT35), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n208_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n282_), .A2(new_n614_), .B1(new_n611_), .B2(new_n610_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n296_), .A2(new_n264_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT73), .B1(new_n616_), .B2(new_n226_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT73), .ZN(new_n618_));
  AOI211_X1 g417(.A(new_n618_), .B(new_n225_), .C1(new_n296_), .C2(new_n264_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n613_), .B(new_n615_), .C1(new_n617_), .C2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n618_), .B1(new_n282_), .B2(new_n225_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n616_), .A2(KEYINPUT73), .A3(new_n226_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n613_), .B1(new_n624_), .B2(new_n615_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n607_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT37), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n615_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n612_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n630_));
  NOR2_X1   g429(.A1(new_n606_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n620_), .A3(new_n631_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n626_), .A2(new_n627_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n627_), .B1(new_n626_), .B2(new_n632_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n603_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n558_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n637_), .A2(G1gat), .A3(new_n556_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT38), .Z(new_n639_));
  NAND2_X1  g438(.A1(new_n516_), .A2(new_n518_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n513_), .A2(new_n514_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n640_), .B(new_n641_), .C1(KEYINPUT33), .C2(new_n481_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n510_), .A2(new_n511_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT98), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n527_), .A2(new_n544_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n547_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n553_), .B1(new_n646_), .B2(new_n453_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n557_), .B1(new_n647_), .B2(new_n383_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n626_), .A2(new_n632_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n648_), .A2(KEYINPUT103), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT103), .B1(new_n648_), .B2(new_n649_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n320_), .A2(KEYINPUT102), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n592_), .A2(new_n594_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n655_), .B(new_n239_), .C1(new_n317_), .C2(new_n319_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n653_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n652_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n527_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G1gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n639_), .A2(new_n660_), .ZN(G1324gat));
  OR3_X1    g460(.A1(new_n637_), .A2(G8gat), .A3(new_n555_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n657_), .B(new_n552_), .C1(new_n651_), .C2(new_n650_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n663_), .A2(new_n664_), .A3(G8gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n663_), .B2(G8gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1325gat));
  INV_X1    g468(.A(new_n637_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n373_), .A3(new_n383_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n658_), .A2(new_n383_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n672_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(new_n672_), .B2(G15gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(G1326gat));
  XOR2_X1   g474(.A(new_n453_), .B(KEYINPUT104), .Z(new_n676_));
  NAND3_X1  g475(.A1(new_n670_), .A2(new_n212_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n658_), .A2(new_n676_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n678_), .A2(G22gat), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n678_), .B2(G22gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(G1327gat));
  AND3_X1   g481(.A1(new_n653_), .A2(new_n656_), .A3(new_n603_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n649_), .A2(KEYINPUT37), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n626_), .A2(new_n627_), .A3(new_n632_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(KEYINPUT106), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n684_), .B1(new_n648_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n635_), .A2(new_n684_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n683_), .B(KEYINPUT44), .C1(new_n691_), .C2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n691_), .A2(new_n693_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n653_), .A2(new_n656_), .A3(new_n603_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(new_n527_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G29gat), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n602_), .A2(new_n649_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n558_), .A2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n556_), .A2(G29gat), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT107), .Z(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n702_), .B2(new_n704_), .ZN(G1328gat));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n694_), .A2(new_n552_), .A3(new_n698_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G36gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n555_), .A2(G36gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n558_), .A2(new_n701_), .A3(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT45), .ZN(new_n713_));
  AOI211_X1 g512(.A(new_n707_), .B(new_n708_), .C1(new_n710_), .C2(new_n713_), .ZN(new_n714_));
  AND4_X1   g513(.A1(KEYINPUT108), .A2(new_n710_), .A3(new_n706_), .A4(new_n713_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  NAND4_X1  g515(.A1(new_n694_), .A2(new_n698_), .A3(G43gat), .A4(new_n383_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n702_), .A2(new_n384_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(G43gat), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g519(.A(new_n676_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n702_), .A2(G50gat), .A3(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n694_), .A2(new_n454_), .A3(new_n698_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(G50gat), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT109), .ZN(G1331gat));
  OR2_X1    g524(.A1(new_n317_), .A2(new_n319_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n239_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n648_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n636_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n527_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n726_), .A2(new_n239_), .A3(new_n603_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n652_), .A2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n556_), .A2(KEYINPUT110), .ZN(new_n735_));
  MUX2_X1   g534(.A(KEYINPUT110), .B(new_n735_), .S(G57gat), .Z(new_n736_));
  AOI21_X1  g535(.A(new_n732_), .B1(new_n734_), .B2(new_n736_), .ZN(G1332gat));
  OAI211_X1 g536(.A(new_n733_), .B(new_n552_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G64gat), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n555_), .A2(G64gat), .ZN(new_n742_));
  OAI22_X1  g541(.A1(new_n740_), .A2(new_n741_), .B1(new_n730_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT111), .ZN(G1333gat));
  NAND3_X1  g543(.A1(new_n731_), .A2(new_n375_), .A3(new_n383_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT49), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n734_), .A2(new_n383_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(G71gat), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT49), .B(new_n375_), .C1(new_n734_), .C2(new_n383_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1334gat));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n734_), .A2(new_n676_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G78gat), .ZN(new_n753_));
  INV_X1    g552(.A(G78gat), .ZN(new_n754_));
  AOI211_X1 g553(.A(KEYINPUT50), .B(new_n754_), .C1(new_n734_), .C2(new_n676_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n676_), .A2(new_n754_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT112), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n753_), .A2(new_n755_), .B1(new_n730_), .B2(new_n757_), .ZN(G1335gat));
  NOR4_X1   g557(.A1(new_n602_), .A2(new_n317_), .A3(new_n319_), .A4(new_n239_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n556_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n729_), .A2(new_n701_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n556_), .A2(G85gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(G1336gat));
  OAI21_X1  g563(.A(G92gat), .B1(new_n760_), .B2(new_n555_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n555_), .A2(G92gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n762_), .B2(new_n766_), .ZN(G1337gat));
  OAI21_X1  g566(.A(G99gat), .B1(new_n760_), .B2(new_n384_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n383_), .A2(new_n249_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n762_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g570(.A1(new_n729_), .A2(new_n250_), .A3(new_n454_), .A4(new_n701_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n454_), .B(new_n759_), .C1(new_n691_), .C2(new_n693_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G106gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G106gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT114), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n772_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n778_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1339gat));
  NOR4_X1   g583(.A1(new_n384_), .A2(new_n556_), .A3(new_n454_), .A4(new_n552_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT119), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT59), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n635_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n239_), .B1(new_n595_), .B2(new_n601_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n319_), .B2(new_n317_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n791_), .B2(KEYINPUT115), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n726_), .B2(new_n790_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT54), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(KEYINPUT115), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n726_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .A4(new_n789_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n795_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n228_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n224_), .A2(new_n227_), .A3(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n205_), .C1(new_n234_), .C2(new_n801_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(new_n235_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n316_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n299_), .B1(new_n304_), .B2(new_n290_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n301_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(KEYINPUT55), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n302_), .A2(new_n809_), .A3(new_n306_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n246_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n245_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT116), .B1(new_n814_), .B2(KEYINPUT56), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n315_), .B(new_n239_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n805_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n649_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n315_), .B(new_n804_), .C1(new_n816_), .C2(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n816_), .A2(new_n825_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n824_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n811_), .A2(new_n246_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n816_), .A2(new_n825_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n315_), .A2(new_n804_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n830_), .A2(KEYINPUT58), .A3(new_n831_), .A4(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n828_), .A2(new_n635_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n823_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT57), .B1(new_n819_), .B2(new_n649_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n603_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n788_), .B1(new_n800_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n786_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n842_));
  AOI211_X1 g641(.A(KEYINPUT116), .B(new_n245_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n825_), .B1(new_n843_), .B2(KEYINPUT117), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n315_), .A2(new_n239_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n817_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n829_), .B2(new_n846_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n844_), .A2(new_n847_), .B1(new_n316_), .B2(new_n804_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n821_), .B1(new_n848_), .B2(new_n820_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n849_), .A2(KEYINPUT118), .A3(new_n823_), .A4(new_n834_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n654_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n842_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n840_), .B1(new_n852_), .B2(new_n800_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n839_), .B(new_n239_), .C1(new_n853_), .C2(new_n787_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G113gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n329_), .A3(new_n239_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1340gat));
  OAI211_X1 g656(.A(new_n839_), .B(new_n727_), .C1(new_n853_), .C2(new_n787_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n327_), .B1(new_n726_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n853_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n327_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1341gat));
  AOI211_X1 g661(.A(new_n603_), .B(new_n840_), .C1(new_n852_), .C2(new_n800_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT120), .B1(new_n863_), .B2(G127gat), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n852_), .A2(new_n800_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n786_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n865_), .B(new_n324_), .C1(new_n867_), .C2(new_n603_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n838_), .B1(new_n867_), .B2(KEYINPUT59), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n851_), .A2(new_n324_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n864_), .A2(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1342gat));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n649_), .B(new_n840_), .C1(new_n852_), .C2(new_n800_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(G134gat), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT121), .B(new_n322_), .C1(new_n867_), .C2(new_n649_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n789_), .A2(new_n322_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n874_), .A2(new_n875_), .B1(new_n869_), .B2(new_n876_), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n383_), .A2(new_n453_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n527_), .A3(new_n555_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT122), .Z(new_n880_));
  NAND2_X1  g679(.A1(new_n866_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n389_), .A3(new_n239_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G141gat), .B1(new_n881_), .B2(new_n728_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n882_), .A2(new_n390_), .A3(new_n727_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G148gat), .B1(new_n881_), .B2(new_n726_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1345gat));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  OR3_X1    g688(.A1(new_n881_), .A2(new_n603_), .A3(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n881_), .B2(new_n603_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1346gat));
  NAND2_X1  g691(.A1(new_n882_), .A2(new_n820_), .ZN(new_n893_));
  INV_X1    g692(.A(G162gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n686_), .B2(new_n689_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n894_), .B1(new_n882_), .B2(new_n895_), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n555_), .A2(new_n527_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n383_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n676_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n728_), .B(new_n900_), .C1(new_n800_), .C2(new_n837_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT22), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(G169gat), .A3(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n354_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1348gat));
  AOI21_X1  g708(.A(new_n900_), .B1(new_n800_), .B2(new_n837_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G176gat), .B1(new_n910_), .B2(new_n727_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n454_), .B1(new_n852_), .B2(new_n800_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n726_), .A2(new_n355_), .A3(new_n898_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1349gat));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n603_), .A2(new_n898_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G183gat), .B1(new_n912_), .B2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n851_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n915_), .B1(new_n917_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n916_), .ZN(new_n922_));
  AOI211_X1 g721(.A(new_n454_), .B(new_n922_), .C1(new_n852_), .C2(new_n800_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n919_), .B(KEYINPUT124), .C1(new_n923_), .C2(G183gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n921_), .A2(new_n924_), .ZN(G1350gat));
  NAND4_X1  g724(.A1(new_n910_), .A2(new_n345_), .A3(new_n347_), .A4(new_n820_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n910_), .A2(new_n635_), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n927_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(KEYINPUT125), .B1(new_n927_), .B2(G190gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n926_), .B1(new_n928_), .B2(new_n929_), .ZN(G1351gat));
  NAND2_X1  g729(.A1(new_n878_), .A2(new_n897_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n852_), .B2(new_n800_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n239_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g733(.A(G204gat), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n932_), .B(new_n727_), .C1(KEYINPUT126), .C2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n932_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n726_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT126), .B(G204gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n936_), .B1(new_n938_), .B2(new_n939_), .ZN(G1353gat));
  NAND2_X1  g739(.A1(new_n932_), .A2(new_n654_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT63), .B(G211gat), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n941_), .B2(new_n944_), .ZN(G1354gat));
  AND3_X1   g744(.A1(new_n932_), .A2(G218gat), .A3(new_n635_), .ZN(new_n946_));
  AOI211_X1 g745(.A(new_n649_), .B(new_n931_), .C1(new_n852_), .C2(new_n800_), .ZN(new_n947_));
  AOI21_X1  g746(.A(G218gat), .B1(new_n947_), .B2(KEYINPUT127), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n949_), .B1(new_n937_), .B2(new_n649_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n946_), .B1(new_n948_), .B2(new_n950_), .ZN(G1355gat));
endmodule


