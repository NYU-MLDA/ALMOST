//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_, new_n969_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n981_, new_n982_, new_n983_, new_n984_, new_n986_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT99), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G169gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(KEYINPUT78), .A2(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(KEYINPUT78), .A2(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT91), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n215_), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(KEYINPUT76), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n214_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(KEYINPUT23), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT92), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n217_), .A2(KEYINPUT76), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n215_), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT23), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n220_), .ZN(new_n228_));
  OAI211_X1 g027(.A(KEYINPUT92), .B(new_n223_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n213_), .B1(new_n224_), .B2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(G197gat), .A2(G204gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT21), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT21), .ZN(new_n235_));
  AND2_X1   g034(.A1(G197gat), .A2(G204gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n234_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT85), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n234_), .A2(new_n238_), .A3(new_n242_), .A4(new_n239_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n239_), .A2(KEYINPUT86), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(new_n234_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(KEYINPUT86), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n241_), .A2(new_n243_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT25), .B(G183gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT89), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT89), .B1(new_n254_), .B2(new_n249_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n248_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n225_), .A2(new_n226_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(KEYINPUT23), .ZN(new_n259_));
  INV_X1    g058(.A(new_n210_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n256_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n231_), .A2(new_n247_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n205_), .B1(new_n266_), .B2(KEYINPUT20), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n241_), .A2(new_n243_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n245_), .A2(new_n246_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n265_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n228_), .B1(new_n258_), .B2(new_n214_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n222_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n212_), .B1(new_n273_), .B2(new_n229_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n205_), .B(KEYINPUT20), .C1(new_n270_), .C2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT26), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n254_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n262_), .B1(new_n279_), .B2(new_n248_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT77), .ZN(new_n281_));
  INV_X1    g080(.A(new_n263_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n281_), .B(new_n282_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n281_), .B1(new_n221_), .B2(new_n282_), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n276_), .A2(new_n277_), .A3(G183gat), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n259_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n209_), .A2(new_n210_), .ZN(new_n288_));
  OAI22_X1  g087(.A1(new_n284_), .A2(new_n285_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n247_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n275_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n204_), .B1(new_n267_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT100), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(KEYINPUT100), .B(new_n204_), .C1(new_n267_), .C2(new_n292_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n204_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT20), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n288_), .B1(new_n259_), .B2(new_n286_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n280_), .A2(new_n283_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT77), .B1(new_n272_), .B2(new_n263_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n298_), .B1(new_n302_), .B2(new_n247_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n259_), .A2(new_n264_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n248_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n252_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n254_), .A2(KEYINPUT89), .A3(new_n249_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT90), .B1(new_n304_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT90), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n256_), .A2(new_n310_), .A3(new_n259_), .A4(new_n264_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT93), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n231_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n274_), .A2(KEYINPUT93), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n297_), .B(new_n303_), .C1(new_n316_), .C2(new_n247_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n295_), .A2(new_n296_), .A3(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G8gat), .B(G36gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT18), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G64gat), .B(G92gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT103), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(KEYINPUT103), .A3(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n303_), .B1(new_n316_), .B2(new_n247_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n204_), .A2(new_n298_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(new_n302_), .B2(new_n247_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n309_), .A2(new_n311_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n273_), .A2(new_n229_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT93), .B1(new_n334_), .B2(new_n213_), .ZN(new_n335_));
  AOI211_X1 g134(.A(new_n313_), .B(new_n212_), .C1(new_n273_), .C2(new_n229_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n247_), .B(new_n333_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT94), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n314_), .A2(new_n315_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(KEYINPUT94), .A3(new_n247_), .A4(new_n333_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n204_), .A2(new_n330_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n329_), .B1(new_n342_), .B2(new_n322_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n328_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n330_), .A2(new_n204_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n337_), .A2(new_n338_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n332_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n323_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n342_), .A2(new_n322_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n329_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT2), .B1(new_n356_), .B2(KEYINPUT82), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT2), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361_));
  INV_X1    g160(.A(G141gat), .ZN(new_n362_));
  INV_X1    g161(.A(G148gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n357_), .A2(new_n360_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n367_), .B1(new_n369_), .B2(KEYINPUT1), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT81), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n374_), .B(new_n367_), .C1(new_n369_), .C2(KEYINPUT1), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT1), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n368_), .A2(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n373_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n356_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n371_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n247_), .B1(KEYINPUT29), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT84), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n386_), .A2(KEYINPUT87), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n386_), .B(KEYINPUT87), .C1(new_n383_), .C2(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n382_), .A2(KEYINPUT29), .ZN(new_n390_));
  XOR2_X1   g189(.A(G22gat), .B(G50gat), .Z(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT83), .B(KEYINPUT28), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n390_), .B(new_n391_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G78gat), .B(G106gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT88), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n389_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n394_), .A2(new_n397_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n399_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n406_), .A2(new_n387_), .A3(new_n388_), .A4(new_n401_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415_));
  INV_X1    g214(.A(G134gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G127gat), .ZN(new_n417_));
  INV_X1    g216(.A(G127gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G134gat), .ZN(new_n419_));
  INV_X1    g218(.A(G120gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G113gat), .ZN(new_n421_));
  INV_X1    g220(.A(G113gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G120gat), .ZN(new_n423_));
  AND4_X1   g222(.A1(new_n417_), .A2(new_n419_), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n417_), .A2(new_n419_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT80), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G127gat), .B(G134gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G113gat), .B(G120gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n372_), .A2(KEYINPUT81), .B1(new_n376_), .B2(new_n368_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n381_), .B1(new_n431_), .B2(new_n375_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n370_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n360_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n357_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n426_), .B(new_n430_), .C1(new_n432_), .C2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n428_), .B(new_n429_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n371_), .B(new_n437_), .C1(new_n378_), .C2(new_n381_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n415_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n430_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n437_), .B2(KEYINPUT80), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT4), .B1(new_n382_), .B2(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n373_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n445_), .A2(new_n380_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n426_), .A2(new_n430_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n424_), .A2(new_n425_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n432_), .A2(new_n435_), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n440_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n414_), .B1(new_n444_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT4), .B1(new_n448_), .B2(new_n450_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n443_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n440_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n413_), .A3(new_n451_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(KEYINPUT101), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT101), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n457_), .A2(new_n460_), .A3(new_n413_), .A4(new_n451_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n442_), .B(KEYINPUT31), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(KEYINPUT79), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465_));
  INV_X1    g264(.A(G15gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT30), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n464_), .B(new_n468_), .Z(new_n469_));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(G43gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n289_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n473_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n408_), .A2(new_n462_), .A3(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n354_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n322_), .A2(KEYINPUT32), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n462_), .B1(new_n318_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n345_), .A2(new_n348_), .A3(new_n479_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT98), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT98), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n345_), .A2(new_n348_), .A3(new_n484_), .A4(new_n479_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n481_), .A2(new_n486_), .A3(KEYINPUT102), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n453_), .A2(KEYINPUT33), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n489_), .B(new_n414_), .C1(new_n444_), .C2(new_n452_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n448_), .A2(new_n450_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n414_), .B1(new_n491_), .B2(new_n456_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n439_), .A2(new_n443_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n456_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT96), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n492_), .B(KEYINPUT96), .C1(new_n493_), .C2(new_n456_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n488_), .A2(new_n490_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT97), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n498_), .A2(new_n350_), .A3(new_n351_), .A4(KEYINPUT97), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n487_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT102), .B1(new_n481_), .B2(new_n486_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n408_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n328_), .A2(new_n343_), .B1(new_n352_), .B2(new_n329_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n462_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n408_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n476_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n478_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT69), .B(G15gat), .ZN(new_n513_));
  INV_X1    g312(.A(G22gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT70), .B(G1gat), .Z(new_n516_));
  INV_X1    g315(.A(G8gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT14), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G1gat), .B(G8gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n518_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n519_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G29gat), .B(G36gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT68), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G43gat), .B(G50gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n524_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n526_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n527_), .A2(new_n531_), .A3(KEYINPUT15), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT15), .B1(new_n527_), .B2(new_n531_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n520_), .B(new_n523_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n523_), .A2(new_n520_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n527_), .A2(new_n531_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n535_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n537_), .A2(new_n523_), .A3(new_n520_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n537_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n535_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G169gat), .B(G197gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n545_), .A2(KEYINPUT73), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT73), .B1(new_n545_), .B2(new_n549_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT74), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n536_), .A2(new_n538_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n541_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n554_), .A2(new_n535_), .B1(new_n534_), .B2(new_n539_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n552_), .B1(new_n555_), .B2(new_n548_), .ZN(new_n556_));
  AND4_X1   g355(.A1(new_n552_), .A2(new_n540_), .A3(new_n544_), .A4(new_n548_), .ZN(new_n557_));
  OAI22_X1  g356(.A1(new_n550_), .A2(new_n551_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n512_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT13), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(KEYINPUT10), .B(G99gat), .Z(new_n563_));
  INV_X1    g362(.A(G106gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G85gat), .B(G92gat), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT9), .ZN(new_n567_));
  INV_X1    g366(.A(G85gat), .ZN(new_n568_));
  INV_X1    g367(.A(G92gat), .ZN(new_n569_));
  OR3_X1    g368(.A1(new_n568_), .A2(new_n569_), .A3(KEYINPUT9), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT6), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n565_), .A2(new_n567_), .A3(new_n570_), .A4(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT7), .ZN(new_n574_));
  AOI211_X1 g373(.A(G99gat), .B(G106gat), .C1(new_n574_), .C2(KEYINPUT65), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(KEYINPUT65), .B2(new_n574_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT64), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n576_), .A2(new_n572_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT8), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n566_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n581_), .B2(new_n566_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n573_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n586_), .A2(KEYINPUT11), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(KEYINPUT11), .ZN(new_n588_));
  XOR2_X1   g387(.A(G71gat), .B(G78gat), .Z(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n585_), .A2(new_n593_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n592_), .B(new_n573_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n562_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT66), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT12), .ZN(new_n599_));
  INV_X1    g398(.A(new_n573_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n581_), .A2(new_n566_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT8), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n581_), .A2(new_n582_), .A3(new_n566_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n600_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n599_), .B1(new_n604_), .B2(new_n592_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT67), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n590_), .A2(new_n606_), .A3(new_n591_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n585_), .A2(new_n610_), .A3(KEYINPUT12), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n605_), .A2(new_n562_), .A3(new_n611_), .A4(new_n595_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n598_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n596_), .A2(new_n597_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT5), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  NOR3_X1   g417(.A1(new_n613_), .A2(new_n614_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n609_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(KEYINPUT12), .A3(new_n607_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n595_), .B1(new_n604_), .B2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT12), .B1(new_n585_), .B2(new_n593_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n625_), .A2(new_n562_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n614_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n620_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n561_), .B1(new_n619_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT34), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n538_), .B(new_n573_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n602_), .A2(new_n603_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT15), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n537_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n527_), .A2(new_n531_), .A3(KEYINPUT15), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n634_), .A2(new_n573_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT35), .B(new_n631_), .C1(new_n633_), .C2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G190gat), .B(G218gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G134gat), .B(G162gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(KEYINPUT36), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n585_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n631_), .A2(KEYINPUT35), .ZN(new_n645_));
  INV_X1    g444(.A(new_n631_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT35), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n644_), .A2(new_n645_), .A3(new_n632_), .A4(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n639_), .A2(new_n643_), .A3(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n642_), .B(KEYINPUT36), .Z(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n639_), .B2(new_n649_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT37), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n639_), .A2(new_n649_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n651_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT37), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n639_), .A2(new_n643_), .A3(new_n649_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT72), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT71), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n523_), .B2(new_n520_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n523_), .A2(new_n662_), .A3(new_n520_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n664_), .A2(G231gat), .A3(G233gat), .A4(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(G231gat), .A2(G233gat), .ZN(new_n667_));
  INV_X1    g466(.A(new_n665_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(new_n663_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n610_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n666_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(G127gat), .B(G155gat), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT16), .ZN(new_n673_));
  XNOR2_X1  g472(.A(G183gat), .B(G211gat), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT17), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n671_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n670_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n661_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n679_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n681_), .A2(KEYINPUT72), .A3(new_n677_), .A4(new_n671_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n666_), .A2(new_n669_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n592_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n666_), .A2(new_n669_), .A3(new_n593_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n675_), .B(KEYINPUT17), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n680_), .A2(new_n682_), .A3(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n618_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n626_), .A2(new_n627_), .A3(new_n620_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(KEYINPUT13), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n629_), .A2(new_n660_), .A3(new_n688_), .A4(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n560_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n507_), .A2(KEYINPUT104), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n507_), .A2(KEYINPUT104), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(new_n516_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT105), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n699_), .A2(KEYINPUT105), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n202_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n702_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT38), .A3(new_n700_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n650_), .A2(new_n653_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT106), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n512_), .A2(new_n708_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n689_), .A2(new_n690_), .A3(KEYINPUT13), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT13), .B1(new_n689_), .B2(new_n690_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n680_), .A2(new_n682_), .A3(new_n687_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n713_), .A2(new_n559_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n709_), .A2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G1gat), .B1(new_n716_), .B2(new_n462_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n703_), .A2(new_n705_), .A3(new_n717_), .ZN(G1324gat));
  NAND3_X1  g517(.A1(new_n695_), .A2(new_n517_), .A3(new_n354_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G8gat), .B1(new_n716_), .B2(new_n506_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT39), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT39), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT40), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT40), .B(new_n719_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1325gat));
  OAI21_X1  g526(.A(G15gat), .B1(new_n716_), .B2(new_n511_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT41), .Z(new_n729_));
  NAND3_X1  g528(.A1(new_n695_), .A2(new_n466_), .A3(new_n476_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1326gat));
  OAI21_X1  g530(.A(G22gat), .B1(new_n716_), .B2(new_n408_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT42), .ZN(new_n733_));
  INV_X1    g532(.A(new_n408_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n514_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT107), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n733_), .B1(new_n694_), .B2(new_n736_), .ZN(G1327gat));
  NAND2_X1  g536(.A1(new_n714_), .A2(new_n706_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT111), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(new_n713_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n560_), .A2(new_n740_), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n741_), .A2(G29gat), .A3(new_n462_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n713_), .A2(new_n559_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n714_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n354_), .A2(new_n477_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n318_), .A2(new_n480_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n484_), .B1(new_n342_), .B2(new_n479_), .ZN(new_n750_));
  AND4_X1   g549(.A1(new_n484_), .A2(new_n345_), .A3(new_n348_), .A4(new_n479_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n749_), .B(new_n507_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT102), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(new_n487_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n755_), .A2(new_n408_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n748_), .B1(new_n756_), .B2(new_n476_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n660_), .B(KEYINPUT108), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n747_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n660_), .A2(KEYINPUT43), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n510_), .A2(new_n511_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n748_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n743_), .B(new_n746_), .C1(new_n759_), .C2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n758_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n512_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n757_), .A2(new_n760_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n745_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n764_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(KEYINPUT110), .A3(new_n698_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G29gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT110), .B1(new_n771_), .B2(new_n698_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n742_), .B1(new_n773_), .B2(new_n774_), .ZN(G1328gat));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n776_));
  INV_X1    g575(.A(G36gat), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n560_), .A2(new_n777_), .A3(new_n354_), .A4(new_n740_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT45), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n777_), .B1(new_n771_), .B2(new_n354_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n776_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n759_), .A2(new_n763_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n769_), .B1(new_n783_), .B2(new_n745_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n506_), .B1(new_n784_), .B2(new_n764_), .ZN(new_n785_));
  OAI211_X1 g584(.A(KEYINPUT46), .B(new_n779_), .C1(new_n785_), .C2(new_n777_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(new_n786_), .ZN(G1329gat));
  INV_X1    g586(.A(G43gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n771_), .B2(new_n476_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n741_), .A2(G43gat), .A3(new_n511_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT47), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n792_));
  INV_X1    g591(.A(new_n790_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n511_), .B1(new_n784_), .B2(new_n764_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n792_), .B(new_n793_), .C1(new_n794_), .C2(new_n788_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1330gat));
  AOI21_X1  g595(.A(new_n408_), .B1(new_n784_), .B2(new_n764_), .ZN(new_n797_));
  INV_X1    g596(.A(G50gat), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n408_), .A2(G50gat), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT112), .ZN(new_n800_));
  OAI22_X1  g599(.A1(new_n797_), .A2(new_n798_), .B1(new_n741_), .B2(new_n800_), .ZN(G1331gat));
  NOR3_X1   g600(.A1(new_n712_), .A2(new_n558_), .A3(new_n714_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n709_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G57gat), .B1(new_n803_), .B2(new_n462_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n512_), .A2(new_n558_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n714_), .B1(new_n659_), .B2(new_n654_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n713_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n698_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n808_), .A2(G57gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n804_), .B1(new_n807_), .B2(new_n809_), .ZN(G1332gat));
  OAI21_X1  g609(.A(G64gat), .B1(new_n803_), .B2(new_n506_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT48), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n506_), .A2(G64gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n807_), .B2(new_n813_), .ZN(G1333gat));
  OAI21_X1  g613(.A(G71gat), .B1(new_n803_), .B2(new_n511_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT49), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n511_), .A2(G71gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n807_), .B2(new_n817_), .ZN(G1334gat));
  OAI21_X1  g617(.A(G78gat), .B1(new_n803_), .B2(new_n408_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT50), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n408_), .A2(G78gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n807_), .B2(new_n821_), .ZN(G1335gat));
  NOR2_X1   g621(.A1(new_n739_), .A2(new_n712_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n805_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n568_), .B1(new_n824_), .B2(new_n808_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT113), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n713_), .A2(new_n559_), .A3(new_n714_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT114), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n783_), .A2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n462_), .A2(new_n568_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n826_), .B1(new_n830_), .B2(new_n831_), .ZN(G1336gat));
  INV_X1    g631(.A(new_n824_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n569_), .A3(new_n354_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n783_), .A2(new_n506_), .A3(new_n829_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n569_), .ZN(G1337gat));
  INV_X1    g635(.A(G99gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n830_), .B2(new_n476_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n833_), .A2(new_n476_), .A3(new_n563_), .ZN(new_n839_));
  OR3_X1    g638(.A1(new_n838_), .A2(new_n839_), .A3(KEYINPUT51), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT51), .B1(new_n838_), .B2(new_n839_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1338gat));
  NAND3_X1  g641(.A1(new_n833_), .A2(new_n564_), .A3(new_n734_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n734_), .B(new_n828_), .C1(new_n759_), .C2(new_n763_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n844_), .A2(new_n845_), .A3(G106gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n844_), .B2(G106gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n843_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g648(.A1(new_n354_), .A2(new_n511_), .A3(new_n808_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n556_), .A2(new_n557_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n534_), .A2(new_n553_), .A3(new_n535_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n554_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n852_), .B(new_n549_), .C1(new_n853_), .C2(new_n535_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n851_), .A2(new_n690_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT55), .B1(new_n562_), .B2(KEYINPUT117), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n562_), .A2(KEYINPUT55), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n605_), .A2(new_n595_), .A3(new_n611_), .A4(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT118), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n858_), .A2(new_n861_), .A3(KEYINPUT118), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT56), .B1(new_n865_), .B2(new_n618_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n858_), .A2(new_n861_), .A3(KEYINPUT118), .ZN(new_n867_));
  OAI211_X1 g666(.A(KEYINPUT56), .B(new_n618_), .C1(new_n867_), .C2(new_n862_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n855_), .B1(new_n866_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n660_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT58), .B(new_n855_), .C1(new_n866_), .C2(new_n869_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n706_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n558_), .A2(new_n690_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n618_), .B1(new_n867_), .B2(new_n862_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT56), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n878_), .B2(new_n868_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n851_), .A2(new_n854_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n874_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n872_), .A2(new_n873_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n874_), .B(KEYINPUT57), .C1(new_n879_), .C2(new_n881_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n688_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n692_), .B2(new_n558_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n693_), .A2(new_n890_), .A3(new_n891_), .A4(new_n559_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n712_), .A2(new_n806_), .A3(new_n891_), .A4(new_n559_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT115), .ZN(new_n894_));
  OAI211_X1 g693(.A(KEYINPUT116), .B(KEYINPUT54), .C1(new_n692_), .C2(new_n558_), .ZN(new_n895_));
  AND4_X1   g694(.A1(new_n889_), .A2(new_n892_), .A3(new_n894_), .A4(new_n895_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n408_), .B(new_n850_), .C1(new_n886_), .C2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(new_n422_), .A3(new_n558_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n870_), .A2(new_n871_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n660_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(new_n904_), .A3(new_n873_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n882_), .A2(new_n883_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(new_n906_), .A3(new_n885_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n714_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n889_), .A2(new_n892_), .A3(new_n894_), .A4(new_n895_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n734_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(KEYINPUT59), .B1(new_n910_), .B2(new_n850_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n900_), .B1(new_n902_), .B2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n897_), .A2(new_n901_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n910_), .A2(KEYINPUT59), .A3(new_n850_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n914_), .A3(KEYINPUT119), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n559_), .B1(new_n912_), .B2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n899_), .B1(new_n916_), .B2(new_n422_), .ZN(G1340gat));
  OAI21_X1  g716(.A(new_n420_), .B1(new_n712_), .B2(KEYINPUT60), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n898_), .B(new_n918_), .C1(KEYINPUT60), .C2(new_n420_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n712_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n420_), .ZN(G1341gat));
  NOR2_X1   g720(.A1(new_n714_), .A2(new_n418_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n912_), .B2(new_n915_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n418_), .B1(new_n897_), .B2(new_n714_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT121), .B1(new_n924_), .B2(new_n927_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n913_), .A2(new_n914_), .A3(KEYINPUT119), .ZN(new_n929_));
  AOI21_X1  g728(.A(KEYINPUT119), .B1(new_n913_), .B2(new_n914_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n922_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n925_), .B(KEYINPUT120), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n928_), .A2(new_n934_), .ZN(G1342gat));
  NAND3_X1  g734(.A1(new_n898_), .A2(new_n416_), .A3(new_n708_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n660_), .B1(new_n912_), .B2(new_n915_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n416_), .ZN(G1343gat));
  NAND2_X1  g737(.A1(new_n908_), .A2(new_n909_), .ZN(new_n939_));
  NOR4_X1   g738(.A1(new_n354_), .A2(new_n408_), .A3(new_n476_), .A4(new_n808_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n558_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n713_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g744(.A1(new_n941_), .A2(new_n688_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT122), .ZN(new_n947_));
  XNOR2_X1  g746(.A(KEYINPUT61), .B(G155gat), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(G1346gat));
  AOI21_X1  g748(.A(G162gat), .B1(new_n941_), .B2(new_n708_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n758_), .A2(G162gat), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n941_), .B2(new_n951_), .ZN(G1347gat));
  INV_X1    g751(.A(new_n910_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n506_), .A2(new_n511_), .A3(new_n698_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(KEYINPUT123), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n953_), .A2(new_n955_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n956_), .A2(new_n206_), .A3(new_n558_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n955_), .A2(new_n559_), .ZN(new_n958_));
  OR2_X1    g757(.A1(new_n958_), .A2(KEYINPUT124), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(KEYINPUT124), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n959_), .A2(new_n910_), .A3(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962_));
  AND3_X1   g761(.A1(new_n961_), .A2(new_n962_), .A3(G169gat), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n962_), .B1(new_n961_), .B2(G169gat), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n957_), .B1(new_n963_), .B2(new_n964_), .ZN(G1348gat));
  NAND2_X1  g764(.A1(new_n956_), .A2(new_n713_), .ZN(new_n966_));
  INV_X1    g765(.A(G176gat), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  AND2_X1   g767(.A1(new_n207_), .A2(new_n208_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(new_n966_), .ZN(G1349gat));
  NAND2_X1  g769(.A1(new_n956_), .A2(new_n688_), .ZN(new_n971_));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n972_), .B2(G183gat), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n248_), .B1(KEYINPUT125), .B2(G183gat), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n971_), .B2(new_n974_), .ZN(G1350gat));
  OAI211_X1 g774(.A(new_n956_), .B(new_n708_), .C1(new_n255_), .C2(new_n253_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n956_), .A2(new_n904_), .ZN(new_n977_));
  AND3_X1   g776(.A1(new_n977_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n978_));
  AOI21_X1  g777(.A(KEYINPUT126), .B1(new_n977_), .B2(G190gat), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n976_), .B1(new_n978_), .B2(new_n979_), .ZN(G1351gat));
  NOR4_X1   g779(.A1(new_n506_), .A2(new_n507_), .A3(new_n408_), .A4(new_n476_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n939_), .A2(new_n981_), .ZN(new_n982_));
  INV_X1    g781(.A(new_n982_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n983_), .A2(new_n558_), .ZN(new_n984_));
  XNOR2_X1  g783(.A(new_n984_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g784(.A1(new_n983_), .A2(new_n713_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n986_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g786(.A(new_n714_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(KEYINPUT127), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n983_), .A2(new_n989_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n991_));
  XOR2_X1   g790(.A(new_n990_), .B(new_n991_), .Z(G1354gat));
  OAI21_X1  g791(.A(G218gat), .B1(new_n982_), .B2(new_n660_), .ZN(new_n993_));
  OR2_X1    g792(.A1(new_n707_), .A2(G218gat), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n993_), .B1(new_n982_), .B2(new_n994_), .ZN(G1355gat));
endmodule


