//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n203_), .B1(KEYINPUT1), .B2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n203_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n219_), .A2(new_n204_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n209_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G211gat), .B(G218gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT87), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G197gat), .B(G204gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT21), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n225_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G197gat), .B(G204gat), .Z(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT21), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n229_), .ZN(new_n235_));
  INV_X1    g034(.A(G218gat), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n236_), .A2(G211gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(G211gat), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT87), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n234_), .B(new_n235_), .C1(new_n226_), .C2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n223_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n223_), .B2(new_n241_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G78gat), .B(G106gat), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n245_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n250_));
  XOR2_X1   g049(.A(G22gat), .B(G50gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT28), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n250_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT88), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n253_), .B1(new_n246_), .B2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n249_), .A2(new_n255_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G1gat), .B(G29gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G85gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G57gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G127gat), .B(G134gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n222_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n265_), .B(new_n266_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n209_), .A3(new_n221_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n270_), .A3(KEYINPUT4), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT94), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G225gat), .A2(G233gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(KEYINPUT93), .B(KEYINPUT4), .Z(new_n275_));
  NAND3_X1  g074(.A1(new_n222_), .A2(new_n267_), .A3(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n271_), .A2(new_n272_), .A3(new_n274_), .A4(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n268_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n274_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n272_), .B1(new_n281_), .B2(new_n271_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n264_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n268_), .A2(KEYINPUT4), .A3(new_n270_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT94), .B1(new_n284_), .B2(new_n280_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n285_), .A2(new_n263_), .A3(new_n278_), .A4(new_n277_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(KEYINPUT97), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT97), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n288_), .B(new_n264_), .C1(new_n279_), .C2(new_n282_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(G183gat), .A3(G190gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n294_), .A2(new_n295_), .A3(KEYINPUT23), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n294_), .B2(KEYINPUT23), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n293_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(KEYINPUT24), .A3(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n299_), .A2(KEYINPUT24), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT25), .B(G183gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT26), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n306_));
  INV_X1    g105(.A(G190gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT26), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n303_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n298_), .A2(new_n301_), .A3(new_n302_), .A4(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n294_), .A2(KEYINPUT23), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n293_), .ZN(new_n312_));
  INV_X1    g111(.A(G183gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n307_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n312_), .A2(new_n314_), .B1(G169gat), .B2(G176gat), .ZN(new_n315_));
  INV_X1    g114(.A(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT22), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT86), .B1(new_n317_), .B2(G169gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT22), .B(G169gat), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n316_), .B(new_n318_), .C1(new_n319_), .C2(KEYINPUT86), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n310_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G71gat), .B(G99gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G43gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n322_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(new_n267_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G227gat), .A2(G233gat), .ZN(new_n327_));
  INV_X1    g126(.A(G15gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT30), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT31), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n326_), .B(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n291_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT27), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n319_), .A2(new_n316_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT90), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n300_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n298_), .A2(KEYINPUT91), .A3(new_n314_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT91), .B1(new_n298_), .B2(new_n314_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n232_), .A2(new_n240_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n303_), .ZN(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT26), .B(G190gat), .Z(new_n345_));
  OAI21_X1  g144(.A(new_n312_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n302_), .A2(new_n301_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n342_), .A2(new_n343_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT20), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n241_), .A2(new_n322_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT20), .B1(new_n241_), .B2(new_n322_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n342_), .A2(new_n349_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n241_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n354_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT92), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n298_), .A2(new_n314_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT91), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n298_), .A2(KEYINPUT91), .A3(new_n314_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n338_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n241_), .B1(new_n366_), .B2(new_n348_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n357_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT92), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(new_n354_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n356_), .B1(new_n361_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT18), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NOR2_X1   g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  AOI211_X1 g177(.A(new_n378_), .B(new_n356_), .C1(new_n361_), .C2(new_n371_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n334_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT96), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n355_), .B1(new_n351_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n350_), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n360_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n369_), .A2(new_n354_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n378_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n372_), .A2(new_n376_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(KEYINPUT27), .ZN(new_n388_));
  AND4_X1   g187(.A1(new_n259_), .A2(new_n333_), .A3(new_n380_), .A4(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n256_), .A2(new_n257_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n380_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT95), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n286_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT33), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n286_), .A2(new_n392_), .A3(KEYINPUT33), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OR3_X1    g196(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n370_), .B1(new_n369_), .B2(new_n354_), .ZN(new_n399_));
  AOI211_X1 g198(.A(KEYINPUT92), .B(new_n360_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n378_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n271_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n268_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n264_), .A3(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n397_), .A2(new_n402_), .A3(new_n387_), .A4(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT32), .B(new_n376_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n376_), .A2(KEYINPUT32), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n372_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n407_), .A2(new_n289_), .A3(new_n409_), .A4(new_n287_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n391_), .B1(new_n411_), .B2(new_n258_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n389_), .B1(new_n412_), .B2(new_n332_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G229gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G15gat), .B(G22gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT80), .B(G8gat), .ZN(new_n417_));
  INV_X1    g216(.A(G1gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G1gat), .B(G8gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n416_), .B(new_n422_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G43gat), .B(G50gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G36gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(G29gat), .ZN(new_n430_));
  INV_X1    g229(.A(G29gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G36gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n432_), .A3(KEYINPUT73), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT73), .B1(new_n430_), .B2(new_n432_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n428_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n432_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT73), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n433_), .A3(new_n427_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n426_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n426_), .A2(new_n442_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n415_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT15), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n436_), .A2(new_n440_), .A3(KEYINPUT15), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n424_), .A2(new_n425_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(new_n443_), .A3(new_n414_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n446_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G113gat), .B(G141gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G169gat), .B(G197gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n446_), .A2(new_n453_), .A3(new_n457_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n461_), .B(KEYINPUT83), .Z(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n202_), .B1(new_n413_), .B2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n380_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n258_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n332_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n380_), .A2(new_n388_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(new_n259_), .A3(new_n333_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT98), .A3(new_n462_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n464_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n307_), .A2(new_n236_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G190gat), .A2(G218gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT75), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT75), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n478_), .A3(new_n475_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G134gat), .B(G162gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n477_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT36), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n479_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n480_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n477_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n483_), .A2(new_n489_), .A3(KEYINPUT77), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT77), .B1(new_n483_), .B2(new_n489_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT78), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT78), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT77), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT36), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n487_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n483_), .A2(new_n489_), .A3(KEYINPUT77), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n493_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n492_), .A2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT6), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT7), .ZN(new_n509_));
  INV_X1    g308(.A(G99gat), .ZN(new_n510_));
  INV_X1    g309(.A(G106gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n503_), .B1(new_n508_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT8), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n517_), .B(new_n503_), .C1(new_n508_), .C2(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n520_));
  AND2_X1   g319(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT65), .B1(new_n523_), .B2(new_n511_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT10), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n510_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n526_), .A2(KEYINPUT65), .A3(new_n511_), .A4(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n524_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(G85gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT9), .ZN(new_n532_));
  AND2_X1   g331(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n501_), .A2(KEYINPUT9), .A3(new_n502_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n505_), .A2(new_n507_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n520_), .B1(new_n530_), .B2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n526_), .A2(new_n511_), .A3(new_n527_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT65), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n528_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(new_n544_), .A3(KEYINPUT67), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n519_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n450_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT35), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n442_), .A2(new_n519_), .A3(new_n539_), .A4(new_n545_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n547_), .A2(KEYINPUT74), .A3(new_n552_), .A4(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT74), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n547_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n551_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n547_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n500_), .B(new_n554_), .C1(new_n557_), .C2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n560_), .A2(KEYINPUT37), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n554_), .B1(new_n559_), .B2(new_n557_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(KEYINPUT76), .A3(new_n495_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT76), .B1(new_n562_), .B2(new_n495_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n561_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(G64gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(G57gat), .ZN(new_n568_));
  INV_X1    g367(.A(G57gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(G64gat), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT68), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n568_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n571_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT11), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n568_), .A2(new_n570_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT68), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT11), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n568_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n574_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(KEYINPUT11), .B(new_n580_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n426_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n583_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n451_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(KEYINPUT81), .A3(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G127gat), .B(G155gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT16), .ZN(new_n593_));
  XOR2_X1   g392(.A(G183gat), .B(G211gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n591_), .B(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n587_), .A2(new_n590_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n596_), .A3(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n562_), .A2(new_n495_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT76), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n562_), .A2(KEYINPUT79), .B1(new_n498_), .B2(new_n497_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT79), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n606_), .B(new_n554_), .C1(new_n559_), .C2(new_n557_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n604_), .A2(new_n563_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n566_), .B(new_n601_), .C1(new_n608_), .C2(KEYINPUT37), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT70), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n546_), .A2(KEYINPUT12), .A3(new_n584_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n540_), .A2(new_n544_), .A3(KEYINPUT67), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT67), .B1(new_n540_), .B2(new_n544_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n588_), .B1(new_n614_), .B2(new_n519_), .ZN(new_n615_));
  XOR2_X1   g414(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n611_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT64), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n546_), .B2(new_n584_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n610_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n546_), .A2(new_n584_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n615_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n546_), .A2(new_n584_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n616_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n626_), .A2(new_n628_), .A3(KEYINPUT70), .A4(new_n611_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n623_), .A2(new_n625_), .A3(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(G120gat), .B(G148gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT72), .ZN(new_n632_));
  XOR2_X1   g431(.A(G176gat), .B(G204gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n630_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT13), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n623_), .A2(new_n625_), .A3(new_n629_), .A4(new_n636_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n609_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT82), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n473_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n418_), .A3(new_n291_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT38), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n461_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n643_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n601_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n608_), .B(KEYINPUT99), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n471_), .A3(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n655_), .B2(new_n290_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n647_), .A2(new_n648_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n649_), .A2(new_n656_), .A3(new_n657_), .ZN(G1324gat));
  NAND4_X1  g457(.A1(new_n473_), .A2(new_n468_), .A3(new_n417_), .A4(new_n645_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n653_), .A2(new_n468_), .A3(new_n471_), .A4(new_n654_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(G8gat), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n660_), .B2(G8gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n659_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT101), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n659_), .B(new_n667_), .C1(new_n664_), .C2(new_n663_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n666_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n655_), .B2(new_n332_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT41), .Z(new_n674_));
  INV_X1    g473(.A(new_n332_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n646_), .A2(new_n328_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1326gat));
  OAI21_X1  g476(.A(G22gat), .B1(new_n655_), .B2(new_n259_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT42), .ZN(new_n679_));
  INV_X1    g478(.A(G22gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n646_), .A2(new_n680_), .A3(new_n258_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT102), .ZN(G1327gat));
  INV_X1    g482(.A(new_n601_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n651_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n651_), .A2(KEYINPUT103), .A3(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n566_), .B1(new_n608_), .B2(KEYINPUT37), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n471_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n691_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT43), .B(new_n693_), .C1(new_n467_), .C2(new_n470_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n689_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT44), .B(new_n689_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n698_));
  AND4_X1   g497(.A1(G29gat), .A2(new_n697_), .A3(new_n291_), .A4(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n684_), .A2(new_n608_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n643_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n473_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G29gat), .B1(new_n702_), .B2(new_n291_), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n699_), .A2(new_n703_), .A3(KEYINPUT104), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT104), .B1(new_n699_), .B2(new_n703_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n468_), .A3(new_n698_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G36gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n469_), .A2(G36gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT98), .B1(new_n471_), .B2(new_n462_), .ZN(new_n710_));
  AOI211_X1 g509(.A(new_n202_), .B(new_n463_), .C1(new_n467_), .C2(new_n470_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n701_), .B(new_n709_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT105), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n473_), .A2(new_n714_), .A3(new_n701_), .A4(new_n709_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n713_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n708_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n708_), .B(KEYINPUT46), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  AND4_X1   g522(.A1(G43gat), .A2(new_n697_), .A3(new_n675_), .A4(new_n698_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT106), .B(G43gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n702_), .B2(new_n675_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n724_), .A2(new_n726_), .A3(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1330gat));
  AOI21_X1  g530(.A(G50gat), .B1(new_n702_), .B2(new_n258_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n697_), .A2(new_n698_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n258_), .A2(G50gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(G1331gat));
  INV_X1    g534(.A(new_n643_), .ZN(new_n736_));
  NOR4_X1   g535(.A1(new_n413_), .A2(new_n461_), .A3(new_n736_), .A4(new_n609_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n569_), .A3(new_n291_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n736_), .A2(new_n462_), .A3(new_n684_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n471_), .A2(new_n654_), .A3(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n290_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n740_), .B2(new_n469_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT48), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n468_), .A2(new_n567_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT108), .Z(new_n746_));
  NAND2_X1  g545(.A1(new_n737_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n747_), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n740_), .B2(new_n332_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT49), .ZN(new_n750_));
  INV_X1    g549(.A(G71gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n737_), .A2(new_n751_), .A3(new_n675_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n740_), .B2(new_n259_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n737_), .A2(new_n756_), .A3(new_n258_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1335gat));
  NOR3_X1   g557(.A1(new_n413_), .A2(new_n461_), .A3(new_n736_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n700_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n531_), .A3(new_n291_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n643_), .A2(new_n650_), .A3(new_n684_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT109), .B1(new_n692_), .B2(new_n694_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n413_), .B2(new_n693_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n471_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n764_), .B1(new_n765_), .B2(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n291_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n763_), .B1(new_n771_), .B2(new_n531_), .ZN(G1336gat));
  AOI21_X1  g571(.A(G92gat), .B1(new_n762_), .B2(new_n468_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n533_), .A2(new_n534_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n469_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n770_), .B2(new_n775_), .ZN(G1337gat));
  AOI21_X1  g575(.A(new_n510_), .B1(new_n770_), .B2(new_n675_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n675_), .A2(new_n523_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n761_), .B2(new_n779_), .ZN(new_n780_));
  OR3_X1    g579(.A1(new_n777_), .A2(KEYINPUT51), .A3(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT51), .B1(new_n777_), .B2(new_n780_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1338gat));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n258_), .A2(new_n511_), .ZN(new_n785_));
  OR3_X1    g584(.A1(new_n761_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n761_), .B2(new_n785_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n764_), .A2(new_n259_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT112), .B1(new_n790_), .B2(new_n511_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n692_), .A2(new_n694_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n792_), .B(G106gat), .C1(new_n793_), .C2(new_n789_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(KEYINPUT52), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT112), .B(new_n796_), .C1(new_n790_), .C2(new_n511_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n788_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT53), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n788_), .A2(new_n795_), .A3(new_n800_), .A4(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1339gat));
  INV_X1    g601(.A(G113gat), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT59), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n644_), .B2(new_n463_), .ZN(new_n806_));
  NOR4_X1   g605(.A1(new_n609_), .A2(new_n643_), .A3(KEYINPUT54), .A4(new_n462_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n414_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n452_), .A2(new_n443_), .A3(new_n415_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n458_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n460_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT113), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n460_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n817_), .A2(new_n640_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n623_), .A2(new_n819_), .A3(new_n629_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n611_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n617_), .B1(new_n546_), .B2(new_n584_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n821_), .A2(new_n622_), .A3(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n614_), .A2(new_n588_), .A3(new_n519_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n628_), .A2(new_n824_), .A3(new_n611_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n823_), .A2(KEYINPUT55), .B1(new_n825_), .B2(new_n620_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n827_), .B2(new_n637_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n829_), .B(new_n636_), .C1(new_n820_), .C2(new_n826_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n818_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n809_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n827_), .A2(new_n637_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n829_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n827_), .A2(KEYINPUT56), .A3(new_n637_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n837_), .A2(KEYINPUT114), .A3(KEYINPUT58), .A4(new_n818_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n831_), .A2(new_n832_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n833_), .A2(new_n838_), .A3(new_n691_), .A4(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n608_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n640_), .A2(new_n461_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n638_), .A2(new_n640_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n817_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n841_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n842_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n845_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT57), .A3(new_n841_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n840_), .A2(new_n849_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n808_), .B1(new_n854_), .B2(new_n684_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n468_), .A2(new_n258_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n291_), .A3(new_n675_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n804_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n857_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(new_n852_), .B2(new_n841_), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n848_), .B(new_n608_), .C1(new_n851_), .C2(new_n845_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n601_), .B1(new_n862_), .B2(new_n840_), .ZN(new_n863_));
  OAI211_X1 g662(.A(KEYINPUT59), .B(new_n859_), .C1(new_n863_), .C2(new_n808_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n858_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n803_), .B1(new_n865_), .B2(new_n462_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n855_), .A2(new_n857_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n461_), .A2(new_n803_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT115), .B1(new_n866_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n463_), .B1(new_n858_), .B2(new_n864_), .ZN(new_n873_));
  OAI221_X1 g672(.A(new_n872_), .B1(new_n868_), .B2(new_n869_), .C1(new_n873_), .C2(new_n803_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(G1340gat));
  XOR2_X1   g674(.A(KEYINPUT116), .B(G120gat), .Z(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n736_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n867_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n876_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n736_), .B1(new_n858_), .B2(new_n864_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n876_), .ZN(G1341gat));
  AOI21_X1  g679(.A(G127gat), .B1(new_n867_), .B2(new_n601_), .ZN(new_n881_));
  INV_X1    g680(.A(G127gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n601_), .B2(KEYINPUT117), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(KEYINPUT117), .B2(new_n882_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n881_), .B1(new_n865_), .B2(new_n884_), .ZN(G1342gat));
  AOI21_X1  g684(.A(new_n693_), .B1(new_n858_), .B2(new_n864_), .ZN(new_n886_));
  INV_X1    g685(.A(G134gat), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n654_), .A2(G134gat), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n886_), .A2(new_n887_), .B1(new_n868_), .B2(new_n888_), .ZN(G1343gat));
  NOR4_X1   g688(.A1(new_n468_), .A2(new_n259_), .A3(new_n290_), .A4(new_n675_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n855_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(new_n893_), .B2(new_n650_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n895_), .A3(new_n461_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT118), .B(G141gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n894_), .A2(new_n896_), .A3(new_n898_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1344gat));
  NAND2_X1  g701(.A1(new_n892_), .A2(new_n643_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT120), .B(G148gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1345gat));
  NAND2_X1  g704(.A1(new_n892_), .A2(new_n601_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT121), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n892_), .A2(new_n908_), .A3(new_n601_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n907_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n893_), .B2(new_n693_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n654_), .A2(G162gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n893_), .B2(new_n915_), .ZN(G1347gat));
  INV_X1    g715(.A(new_n855_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n468_), .A2(new_n333_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n650_), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT122), .Z(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(new_n259_), .A3(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n921_), .A2(new_n922_), .A3(G169gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n921_), .B2(G169gat), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n918_), .A2(new_n258_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT123), .B1(new_n855_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n855_), .A2(KEYINPUT123), .A3(new_n927_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n461_), .A2(new_n319_), .ZN(new_n932_));
  OAI22_X1  g731(.A1(new_n924_), .A2(new_n925_), .B1(new_n931_), .B2(new_n932_), .ZN(G1348gat));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n855_), .A2(new_n927_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n316_), .B1(new_n935_), .B2(new_n643_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n736_), .A2(G176gat), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n934_), .B(new_n937_), .C1(new_n931_), .C2(new_n939_), .ZN(new_n940_));
  OR3_X1    g739(.A1(new_n855_), .A2(KEYINPUT123), .A3(new_n927_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n939_), .B1(new_n941_), .B2(new_n928_), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT124), .B1(new_n942_), .B2(new_n936_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n940_), .A2(new_n943_), .ZN(G1349gat));
  AOI211_X1 g743(.A(new_n303_), .B(new_n684_), .C1(new_n941_), .C2(new_n928_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n935_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n946_), .A2(KEYINPUT125), .A3(new_n684_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(G183gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(KEYINPUT125), .B1(new_n946_), .B2(new_n684_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n945_), .B1(new_n948_), .B2(new_n949_), .ZN(G1350gat));
  OAI21_X1  g749(.A(G190gat), .B1(new_n931_), .B2(new_n693_), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n654_), .A2(new_n345_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n931_), .B2(new_n952_), .ZN(G1351gat));
  NAND3_X1  g752(.A1(new_n468_), .A2(new_n390_), .A3(new_n332_), .ZN(new_n954_));
  OR3_X1    g753(.A1(new_n855_), .A2(KEYINPUT126), .A3(new_n954_), .ZN(new_n955_));
  OAI21_X1  g754(.A(KEYINPUT126), .B1(new_n855_), .B2(new_n954_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n955_), .A2(new_n956_), .ZN(new_n957_));
  AND3_X1   g756(.A1(new_n957_), .A2(G197gat), .A3(new_n461_), .ZN(new_n958_));
  AOI21_X1  g757(.A(G197gat), .B1(new_n957_), .B2(new_n461_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1352gat));
  INV_X1    g759(.A(new_n957_), .ZN(new_n961_));
  OAI21_X1  g760(.A(G204gat), .B1(new_n961_), .B2(new_n736_), .ZN(new_n962_));
  INV_X1    g761(.A(G204gat), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n957_), .A2(new_n963_), .A3(new_n643_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(G1353gat));
  AOI21_X1  g764(.A(new_n684_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(KEYINPUT127), .ZN(new_n968_));
  AND3_X1   g767(.A1(new_n957_), .A2(new_n966_), .A3(new_n968_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(new_n957_), .B2(new_n966_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1354gat));
  OR2_X1    g770(.A1(new_n654_), .A2(G218gat), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n693_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n973_));
  OAI22_X1  g772(.A1(new_n961_), .A2(new_n972_), .B1(new_n973_), .B2(new_n236_), .ZN(G1355gat));
endmodule


