//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n205_), .A2(KEYINPUT78), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(KEYINPUT78), .ZN(new_n207_));
  OAI21_X1  g006(.A(G183gat), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT79), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n210_), .B(G183gat), .C1(new_n206_), .C2(new_n207_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n205_), .A2(G183gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT80), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n209_), .A2(KEYINPUT80), .A3(new_n211_), .A4(new_n214_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT81), .B(KEYINPUT23), .Z(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(new_n219_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G169gat), .B(G176gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(new_n223_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n217_), .A2(new_n218_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n219_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT23), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(new_n221_), .B2(new_n231_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(G183gat), .B2(G190gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n235_));
  OR3_X1    g034(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G99gat), .ZN(new_n238_));
  INV_X1    g037(.A(G43gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n230_), .A2(new_n237_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n241_), .B1(new_n230_), .B2(new_n237_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246_));
  INV_X1    g045(.A(G15gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT30), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT82), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT31), .ZN(new_n252_));
  INV_X1    g051(.A(new_n250_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n252_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n204_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n204_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(new_n255_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT3), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT2), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n263_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n265_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n268_), .B1(new_n269_), .B2(KEYINPUT1), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n273_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n260_), .B1(new_n271_), .B2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n276_), .A2(new_n278_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n281_), .B(new_n204_), .C1(new_n282_), .C2(new_n273_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT93), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n290_), .B(new_n260_), .C1(new_n271_), .C2(new_n279_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n287_), .B(new_n291_), .C1(new_n284_), .C2(new_n290_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G29gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(G85gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT0), .B(G57gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  NAND3_X1  g095(.A1(new_n289_), .A2(new_n292_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT96), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n289_), .A2(new_n292_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n296_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT96), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n289_), .A2(new_n292_), .A3(new_n302_), .A4(new_n296_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n262_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G197gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G204gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n306_), .A2(G204gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT21), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT84), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n306_), .B2(G204gat), .ZN(new_n312_));
  INV_X1    g111(.A(G204gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT84), .A3(G197gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(new_n314_), .A3(new_n307_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT85), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n316_), .A2(new_n317_), .ZN(new_n319_));
  OAI221_X1 g118(.A(new_n310_), .B1(KEYINPUT21), .B2(new_n315_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n316_), .B(KEYINPUT85), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(KEYINPUT21), .A3(new_n315_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n230_), .A2(new_n323_), .A3(new_n237_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n212_), .A2(KEYINPUT89), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n212_), .A2(KEYINPUT89), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT25), .B(G183gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n227_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n233_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n236_), .A2(new_n235_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT91), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n222_), .A2(new_n337_), .ZN(new_n338_));
  OAI22_X1  g137(.A1(new_n329_), .A2(new_n333_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT92), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n320_), .A2(new_n322_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT20), .B(new_n324_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  AOI21_X1  g151(.A(new_n323_), .B1(new_n230_), .B2(new_n237_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT20), .B1(new_n339_), .B2(new_n341_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n347_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n348_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n347_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n358_));
  OAI211_X1 g157(.A(KEYINPUT95), .B(new_n358_), .C1(new_n345_), .C2(new_n347_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(KEYINPUT95), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(KEYINPUT27), .B(new_n357_), .C1(new_n361_), .C2(new_n352_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT27), .ZN(new_n363_));
  INV_X1    g162(.A(new_n347_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT20), .ZN(new_n365_));
  INV_X1    g164(.A(new_n333_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n222_), .A2(new_n337_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n334_), .B(KEYINPUT91), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n366_), .A2(new_n328_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT92), .B1(new_n369_), .B2(new_n323_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n365_), .B1(new_n370_), .B2(new_n342_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n364_), .B1(new_n371_), .B2(new_n324_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n352_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n355_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n352_), .B1(new_n348_), .B2(new_n356_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n363_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n362_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT29), .B1(new_n271_), .B2(new_n279_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n341_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n381_), .A3(new_n341_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G78gat), .B(G106gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n383_), .A2(new_n384_), .A3(KEYINPUT87), .A4(new_n386_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n379_), .A2(new_n381_), .A3(new_n341_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n381_), .B1(new_n379_), .B2(new_n341_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT86), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n383_), .A2(new_n384_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n397_), .A3(new_n385_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n271_), .A2(new_n279_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT28), .ZN(new_n402_));
  NOR4_X1   g201(.A1(new_n271_), .A2(new_n279_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G22gat), .B(G50gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT28), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n409_), .B2(new_n403_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n398_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT88), .B1(new_n392_), .B2(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n398_), .A2(new_n411_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT88), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n391_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n383_), .A2(new_n384_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n385_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n387_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n411_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n413_), .A2(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n305_), .A2(new_n378_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n419_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n415_), .B1(new_n414_), .B2(new_n391_), .ZN(new_n424_));
  AND4_X1   g223(.A1(new_n415_), .A2(new_n391_), .A3(new_n411_), .A4(new_n398_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n377_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n413_), .A2(new_n416_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n348_), .A2(new_n356_), .A3(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n304_), .B(new_n430_), .C1(new_n361_), .C2(new_n429_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n297_), .B(KEYINPUT33), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n373_), .B1(new_n372_), .B2(new_n355_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n296_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT94), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n288_), .B(new_n291_), .C1(new_n284_), .C2(new_n290_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n435_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n432_), .A2(new_n433_), .A3(new_n439_), .A4(new_n357_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n428_), .A2(new_n431_), .A3(new_n440_), .A4(new_n423_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n427_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n304_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n262_), .B1(new_n421_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n422_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT71), .B(G1gat), .ZN(new_n446_));
  INV_X1    g245(.A(G8gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT14), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G15gat), .B(G22gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT72), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT72), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(new_n452_), .A3(new_n449_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G1gat), .B(G8gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n451_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G29gat), .B(G36gat), .Z(new_n459_));
  XOR2_X1   g258(.A(G43gat), .B(G50gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT15), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n457_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n455_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n461_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT77), .ZN(new_n469_));
  OR3_X1    g268(.A1(new_n456_), .A2(new_n461_), .A3(new_n457_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n467_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  AOI211_X1 g272(.A(KEYINPUT77), .B(new_n467_), .C1(new_n466_), .C2(new_n470_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n468_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G113gat), .B(G141gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G169gat), .B(G197gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n468_), .B(new_n478_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n445_), .A2(KEYINPUT97), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT97), .B1(new_n445_), .B2(new_n482_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G230gat), .A2(G233gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT64), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(G85gat), .A2(G92gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT6), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(G99gat), .A3(G106gat), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n497_));
  INV_X1    g296(.A(G99gat), .ZN(new_n498_));
  INV_X1    g297(.A(G106gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n491_), .B1(new_n496_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT8), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n493_), .A2(new_n495_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(new_n501_), .A3(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT8), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n491_), .ZN(new_n508_));
  OR2_X1    g307(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n499_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(KEYINPUT65), .A3(new_n499_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n489_), .A2(KEYINPUT9), .A3(new_n490_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n490_), .A2(KEYINPUT9), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n519_), .A2(new_n505_), .A3(new_n520_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n504_), .A2(new_n508_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT66), .B(G71gat), .ZN(new_n523_));
  INV_X1    g322(.A(G78gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(G71gat), .ZN(new_n527_));
  INV_X1    g326(.A(G71gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(KEYINPUT66), .ZN(new_n529_));
  OAI21_X1  g328(.A(G78gat), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G64gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(G57gat), .ZN(new_n533_));
  INV_X1    g332(.A(G57gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(G64gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n535_), .A3(KEYINPUT11), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT11), .B1(new_n533_), .B2(new_n535_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n530_), .B(new_n525_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n522_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n522_), .A2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n488_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT12), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n518_), .A2(new_n521_), .A3(KEYINPUT67), .ZN(new_n548_));
  INV_X1    g347(.A(new_n508_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n507_), .B1(new_n506_), .B2(new_n491_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT67), .B1(new_n518_), .B2(new_n521_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n547_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n546_), .B1(new_n522_), .B2(new_n541_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n487_), .A4(new_n542_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n545_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G120gat), .B(G148gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n545_), .A2(new_n555_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT69), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n566_), .A2(KEYINPUT69), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n565_), .B1(new_n569_), .B2(new_n567_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n518_), .A2(new_n521_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT67), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n504_), .A2(new_n508_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n548_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n462_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n578_), .A2(KEYINPUT70), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n462_), .A2(new_n577_), .B1(new_n461_), .B2(new_n522_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT34), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n583_));
  OR3_X1    g382(.A1(new_n579_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n580_), .B(new_n585_), .C1(new_n579_), .C2(new_n583_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n590_), .A2(new_n591_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n584_), .A2(new_n591_), .A3(new_n590_), .A4(new_n586_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT37), .B1(new_n594_), .B2(new_n595_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT73), .Z(new_n602_));
  AND2_X1   g401(.A1(new_n465_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n465_), .A2(new_n602_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n541_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n541_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT75), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n613_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT17), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n609_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n616_), .B(new_n617_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n608_), .A3(new_n607_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n600_), .A2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT76), .Z(new_n624_));
  NOR3_X1   g423(.A1(new_n485_), .A2(new_n572_), .A3(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n304_), .A2(new_n446_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n445_), .A2(new_n596_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n571_), .A2(new_n482_), .A3(new_n622_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT98), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT99), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n634_), .B2(new_n443_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n625_), .A2(KEYINPUT38), .A3(new_n626_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n629_), .A2(new_n635_), .A3(new_n636_), .ZN(G1324gat));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n377_), .A3(new_n632_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G8gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT39), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n625_), .A2(new_n447_), .A3(new_n377_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1325gat));
  OAI21_X1  g443(.A(G15gat), .B1(new_n634_), .B2(new_n262_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n262_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n625_), .A2(new_n247_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1326gat));
  OAI21_X1  g449(.A(G22gat), .B1(new_n634_), .B2(new_n421_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n625_), .A2(new_n653_), .A3(new_n426_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1327gat));
  INV_X1    g454(.A(new_n596_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n622_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n485_), .A2(new_n572_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G29gat), .B1(new_n659_), .B2(new_n304_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  INV_X1    g460(.A(new_n600_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n445_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT102), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n445_), .A2(new_n665_), .A3(new_n661_), .A4(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n445_), .A2(new_n662_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n657_), .A2(new_n482_), .A3(new_n571_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT101), .Z(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT44), .B1(new_n669_), .B2(new_n671_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n304_), .A2(G29gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n660_), .B1(new_n674_), .B2(new_n675_), .ZN(G1328gat));
  NOR2_X1   g475(.A1(new_n658_), .A2(new_n572_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n377_), .A2(KEYINPUT103), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n377_), .A2(KEYINPUT103), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(G36gat), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n677_), .B(new_n682_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT45), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n672_), .A2(new_n673_), .A3(new_n378_), .ZN(new_n685_));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT46), .B(new_n684_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1329gat));
  NOR4_X1   g490(.A1(new_n672_), .A2(new_n673_), .A3(new_n239_), .A4(new_n262_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G43gat), .B1(new_n659_), .B2(new_n648_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT47), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n674_), .A2(G43gat), .A3(new_n648_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n693_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n698_), .ZN(G1330gat));
  AOI21_X1  g498(.A(G50gat), .B1(new_n659_), .B2(new_n426_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n426_), .A2(G50gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n674_), .B2(new_n701_), .ZN(G1331gat));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n480_), .A2(new_n481_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n445_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n445_), .B2(new_n704_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n707_), .A2(new_n571_), .A3(new_n624_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n534_), .A3(new_n304_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n630_), .A2(new_n704_), .A3(new_n572_), .A4(new_n622_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n443_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1332gat));
  OAI21_X1  g511(.A(G64gat), .B1(new_n710_), .B2(new_n681_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT48), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n708_), .A2(new_n532_), .A3(new_n680_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1333gat));
  OAI21_X1  g515(.A(G71gat), .B1(new_n710_), .B2(new_n262_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT49), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n708_), .A2(new_n528_), .A3(new_n648_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1334gat));
  OAI21_X1  g519(.A(G78gat), .B1(new_n710_), .B2(new_n421_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n426_), .A2(new_n524_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT106), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n708_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1335gat));
  NOR3_X1   g526(.A1(new_n571_), .A2(new_n482_), .A3(new_n622_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n669_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(G85gat), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n443_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n658_), .A2(new_n571_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n732_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT107), .B(new_n732_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G85gat), .B1(new_n737_), .B2(new_n304_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT108), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT108), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n731_), .B1(new_n739_), .B2(new_n740_), .ZN(G1336gat));
  OAI21_X1  g540(.A(G92gat), .B1(new_n729_), .B2(new_n681_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n737_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n378_), .A2(G92gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n742_), .B1(new_n743_), .B2(new_n744_), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n729_), .B2(new_n262_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n648_), .A2(new_n516_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n737_), .B2(new_n749_), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT109), .B(new_n748_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n746_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT51), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n746_), .B(new_n754_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1338gat));
  XNOR2_X1  g555(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n669_), .A2(new_n426_), .A3(new_n728_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G106gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n760_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(G106gat), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n737_), .A2(new_n499_), .A3(new_n426_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n757_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n758_), .A2(G106gat), .A3(new_n762_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n762_), .B1(new_n758_), .B2(G106gat), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n765_), .B(new_n757_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n766_), .A2(new_n770_), .ZN(G1339gat));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n622_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n572_), .B2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n704_), .A2(KEYINPUT112), .A3(new_n571_), .A4(new_n622_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n600_), .A3(new_n775_), .ZN(new_n776_));
  OR2_X1    g575(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT114), .Z(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n777_), .A3(new_n780_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n471_), .A2(new_n467_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n463_), .A2(new_n466_), .A3(new_n472_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n479_), .A3(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n481_), .A2(new_n564_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n555_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n553_), .A2(new_n554_), .A3(new_n542_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n488_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n577_), .A2(new_n547_), .B1(new_n522_), .B2(new_n541_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n793_), .A2(KEYINPUT55), .A3(new_n487_), .A4(new_n554_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n790_), .A2(new_n792_), .A3(new_n794_), .A4(KEYINPUT115), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n561_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n563_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT56), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n788_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT58), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n788_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n803_), .A2(KEYINPUT56), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n801_), .B(new_n563_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(KEYINPUT117), .A3(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n807_), .A2(new_n662_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n481_), .A2(new_n565_), .A3(new_n787_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n800_), .A2(KEYINPUT116), .A3(new_n801_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n803_), .B2(KEYINPUT56), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n804_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n482_), .A2(new_n564_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n818_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n817_), .B1(new_n825_), .B2(new_n656_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n822_), .A2(new_n824_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT57), .B(new_n596_), .C1(new_n827_), .C2(new_n818_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n807_), .A2(new_n662_), .A3(KEYINPUT118), .A4(new_n813_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n816_), .A2(new_n826_), .A3(new_n828_), .A4(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n784_), .B1(new_n830_), .B2(new_n657_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n426_), .A2(new_n377_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n262_), .A2(new_n443_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT59), .B1(new_n831_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n828_), .A2(new_n826_), .A3(new_n814_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n657_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n782_), .A2(new_n783_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n834_), .A2(KEYINPUT59), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n835_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842_), .B2(new_n704_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n831_), .A2(new_n834_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n704_), .A2(G113gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n843_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  NAND3_X1  g646(.A1(new_n835_), .A2(new_n572_), .A3(new_n841_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT119), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n835_), .A2(new_n850_), .A3(new_n841_), .A4(new_n572_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(G120gat), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(G120gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n571_), .B2(KEYINPUT60), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n844_), .B(new_n854_), .C1(KEYINPUT60), .C2(new_n853_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n855_), .ZN(G1341gat));
  OAI21_X1  g655(.A(G127gat), .B1(new_n842_), .B2(new_n657_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n657_), .A2(G127gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n845_), .B2(new_n858_), .ZN(G1342gat));
  OAI21_X1  g658(.A(G134gat), .B1(new_n842_), .B2(new_n600_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n596_), .A2(G134gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n845_), .B2(new_n861_), .ZN(G1343gat));
  NAND2_X1  g661(.A1(new_n830_), .A2(new_n657_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n838_), .ZN(new_n864_));
  NOR4_X1   g663(.A1(new_n680_), .A2(new_n421_), .A3(new_n443_), .A4(new_n648_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n704_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT120), .B(G141gat), .Z(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1344gat));
  INV_X1    g668(.A(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n572_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n866_), .A2(new_n657_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT61), .B(G155gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  OR3_X1    g674(.A1(new_n866_), .A2(G162gat), .A3(new_n596_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G162gat), .B1(new_n866_), .B2(new_n600_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1347gat));
  NAND2_X1  g677(.A1(new_n680_), .A2(new_n305_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n839_), .A2(new_n482_), .A3(new_n421_), .A4(new_n880_), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT22), .B(G169gat), .Z(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n881_), .B2(G169gat), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n883_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n885_), .A2(new_n886_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n881_), .A2(new_n884_), .A3(G169gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(G1348gat));
  NAND2_X1  g689(.A1(new_n839_), .A2(new_n421_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n879_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G176gat), .B1(new_n892_), .B2(new_n572_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n829_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n811_), .A2(KEYINPUT117), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n600_), .B1(new_n895_), .B2(KEYINPUT58), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT118), .B1(new_n896_), .B2(new_n813_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n894_), .A2(new_n897_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n828_), .A2(new_n826_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n622_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT122), .B(new_n421_), .C1(new_n900_), .C2(new_n784_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n831_), .B2(new_n426_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n879_), .A2(new_n225_), .A3(new_n571_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n893_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  NOR2_X1   g705(.A1(new_n879_), .A2(new_n657_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n891_), .A2(new_n327_), .A3(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n901_), .B2(new_n903_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911_));
  AOI21_X1  g710(.A(G183gat), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(KEYINPUT122), .B1(new_n864_), .B2(new_n421_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n831_), .A2(new_n902_), .A3(new_n426_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n907_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT123), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n909_), .B1(new_n912_), .B2(new_n916_), .ZN(G1350gat));
  AND3_X1   g716(.A1(new_n656_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n839_), .A2(new_n421_), .A3(new_n880_), .A4(new_n918_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n891_), .A2(new_n600_), .A3(new_n879_), .ZN(new_n920_));
  INV_X1    g719(.A(G190gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT124), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n924_), .B(new_n919_), .C1(new_n920_), .C2(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1351gat));
  NOR3_X1   g725(.A1(new_n648_), .A2(new_n421_), .A3(new_n304_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n928_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n929_), .A2(new_n681_), .A3(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n864_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n704_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n306_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n571_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n313_), .ZN(G1353gat));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n864_), .A2(new_n931_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n622_), .ZN(new_n939_));
  XOR2_X1   g738(.A(KEYINPUT63), .B(G211gat), .Z(new_n940_));
  NOR3_X1   g739(.A1(new_n932_), .A2(new_n657_), .A3(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(KEYINPUT126), .B1(new_n939_), .B2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n940_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n938_), .A2(new_n622_), .A3(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n932_), .A2(new_n657_), .ZN(new_n946_));
  OAI211_X1 g745(.A(new_n944_), .B(new_n945_), .C1(new_n946_), .C2(new_n937_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n942_), .A2(new_n947_), .ZN(G1354gat));
  INV_X1    g747(.A(G218gat), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n949_), .B1(new_n938_), .B2(new_n662_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n656_), .A2(new_n949_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n932_), .A2(new_n951_), .ZN(new_n952_));
  OAI21_X1  g751(.A(KEYINPUT127), .B1(new_n950_), .B2(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G218gat), .B1(new_n932_), .B2(new_n600_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955_));
  OAI211_X1 g754(.A(new_n954_), .B(new_n955_), .C1(new_n932_), .C2(new_n951_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n953_), .A2(new_n956_), .ZN(G1355gat));
endmodule


