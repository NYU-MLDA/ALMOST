//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT74), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G134gat), .ZN(new_n204_));
  INV_X1    g003(.A(G162gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT36), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G232gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT72), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT34), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT35), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  OAI21_X1  g017(.A(new_n217_), .B1(new_n218_), .B2(new_n214_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT64), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT10), .B(G99gat), .Z(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  AOI211_X1 g023(.A(new_n221_), .B(new_n222_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n226_), .B(new_n217_), .C1(new_n218_), .C2(new_n214_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n222_), .A2(new_n221_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n224_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n234_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n218_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n241_), .B2(new_n218_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT8), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT67), .B(KEYINPUT8), .Z(new_n247_));
  NAND3_X1  g046(.A1(new_n241_), .A2(new_n218_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n228_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G29gat), .B(G36gat), .Z(new_n251_));
  XOR2_X1   g050(.A(G43gat), .B(G50gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT15), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n213_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n212_), .A2(KEYINPUT35), .ZN(new_n256_));
  INV_X1    g055(.A(new_n228_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n241_), .A2(new_n218_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT68), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n241_), .A2(new_n242_), .A3(new_n218_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT8), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n257_), .B1(new_n261_), .B2(new_n248_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT73), .B1(new_n262_), .B2(new_n253_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n245_), .B1(new_n258_), .B2(KEYINPUT68), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n249_), .B1(new_n264_), .B2(new_n260_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n266_));
  INV_X1    g065(.A(new_n253_), .ZN(new_n267_));
  NOR4_X1   g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n257_), .A4(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n255_), .B(new_n256_), .C1(new_n263_), .C2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n228_), .B(new_n253_), .C1(new_n246_), .C2(new_n249_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n266_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n262_), .A2(KEYINPUT73), .A3(new_n253_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n256_), .B1(new_n274_), .B2(new_n255_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n209_), .B1(new_n270_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n255_), .B1(new_n263_), .B2(new_n268_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n256_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n279_), .A2(new_n207_), .A3(new_n206_), .A4(new_n269_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT105), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(G155gat), .B2(G162gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT3), .Z(new_n289_));
  NAND2_X1  g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(KEYINPUT2), .Z(new_n291_));
  OAI21_X1  g090(.A(new_n287_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n288_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT1), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n290_), .B(new_n293_), .C1(new_n286_), .C2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT86), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G127gat), .B(G134gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G113gat), .B(G120gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT83), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n299_), .B(new_n300_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(KEYINPUT83), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n305_), .A2(KEYINPUT4), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n292_), .A2(new_n296_), .A3(new_n303_), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT96), .Z(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT4), .B1(new_n305_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n306_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n305_), .A2(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n307_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT0), .ZN(new_n317_));
  INV_X1    g116(.A(G57gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(new_n215_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n312_), .A2(new_n320_), .A3(new_n314_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G183gat), .ZN(new_n326_));
  INV_X1    g125(.A(G190gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT23), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT80), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OR3_X1    g129(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT23), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n329_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n327_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT22), .B(G169gat), .ZN(new_n337_));
  INV_X1    g136(.A(G176gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT25), .B(G183gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT26), .B(G190gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(KEYINPUT24), .A3(new_n336_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n344_), .A2(KEYINPUT24), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n343_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n331_), .A2(new_n328_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n340_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G197gat), .B(G204gat), .Z(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT21), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G197gat), .B(G204gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT21), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G211gat), .B(G218gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(KEYINPUT90), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n352_), .A2(new_n356_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(KEYINPUT90), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n350_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(KEYINPUT91), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n347_), .A2(new_n333_), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n339_), .B(KEYINPUT81), .Z(new_n365_));
  NAND2_X1  g164(.A1(new_n348_), .A2(new_n334_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n336_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n364_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(KEYINPUT20), .B(new_n362_), .C1(new_n363_), .C2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT19), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G64gat), .B(G92gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n363_), .A2(new_n368_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n350_), .A2(new_n361_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(new_n371_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(KEYINPUT20), .A3(new_n380_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n372_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n361_), .B(KEYINPUT93), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n350_), .B(KEYINPUT101), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n378_), .B(KEYINPUT20), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n371_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT102), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(KEYINPUT102), .A3(new_n371_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n369_), .A2(new_n371_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n390_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT103), .B(new_n384_), .C1(new_n394_), .C2(new_n377_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT103), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n392_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n377_), .B1(new_n397_), .B2(new_n391_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n382_), .A2(new_n383_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n396_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n372_), .A2(new_n381_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(new_n377_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n402_), .A2(KEYINPUT27), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n395_), .A2(new_n400_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT89), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n297_), .B(new_n408_), .ZN(new_n409_));
  OAI221_X1 g208(.A(new_n363_), .B1(new_n406_), .B2(new_n405_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n411_));
  NAND2_X1  g210(.A1(new_n297_), .A2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n385_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n405_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n410_), .A2(new_n406_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT94), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT28), .B1(new_n298_), .B2(KEYINPUT29), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT28), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n409_), .A2(new_n424_), .A3(new_n407_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT87), .ZN(new_n427_));
  XOR2_X1   g226(.A(G22gat), .B(G50gat), .Z(new_n428_));
  INV_X1    g227(.A(KEYINPUT87), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n423_), .A2(new_n429_), .A3(new_n425_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n428_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n427_), .A2(new_n430_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n428_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT88), .B1(new_n438_), .B2(new_n431_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n422_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n417_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n419_), .A2(new_n431_), .A3(new_n438_), .A4(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n368_), .B(KEYINPUT82), .ZN(new_n443_));
  XOR2_X1   g242(.A(G71gat), .B(G99gat), .Z(new_n444_));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n443_), .B(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G15gat), .B(G43gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT30), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n304_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n449_), .B(new_n453_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n440_), .A2(new_n442_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n325_), .B(new_n404_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n320_), .B1(new_n313_), .B2(new_n307_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT97), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT97), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n460_), .B(new_n320_), .C1(new_n313_), .C2(new_n307_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n308_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT98), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n459_), .B(new_n461_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n462_), .A2(new_n463_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n402_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n320_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT33), .ZN(new_n468_));
  INV_X1    g267(.A(new_n401_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n377_), .A2(KEYINPUT32), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n470_), .B(KEYINPUT99), .Z(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(KEYINPUT100), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n471_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT100), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n324_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n394_), .A2(new_n470_), .ZN(new_n477_));
  OAI22_X1  g276(.A1(new_n466_), .A2(new_n468_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n440_), .A2(new_n442_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n454_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n283_), .B1(new_n457_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT70), .ZN(new_n484_));
  XOR2_X1   g283(.A(G57gat), .B(G64gat), .Z(new_n485_));
  INV_X1    g284(.A(KEYINPUT11), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G57gat), .B(G64gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G71gat), .B(G78gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(new_n490_), .A3(KEYINPUT11), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n492_), .A2(KEYINPUT69), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT69), .B1(new_n492_), .B2(new_n493_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n484_), .B1(new_n250_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n496_), .B1(new_n265_), .B2(new_n257_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n494_), .A2(new_n495_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n262_), .A2(KEYINPUT70), .A3(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(G230gat), .A2(G233gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n262_), .B2(new_n499_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n502_), .B1(new_n262_), .B2(new_n499_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n492_), .A2(new_n493_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(new_n504_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n250_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G120gat), .B(G148gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT71), .B(G204gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT5), .B(G176gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n516_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n503_), .A2(new_n510_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT13), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(KEYINPUT13), .A3(new_n519_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525_));
  INV_X1    g324(.A(G1gat), .ZN(new_n526_));
  INV_X1    g325(.A(G8gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G1gat), .B(G8gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n254_), .A2(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n267_), .A2(new_n531_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n267_), .B(new_n531_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(G197gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT78), .B(G169gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(KEYINPUT77), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n539_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n524_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n531_), .B(new_n548_), .Z(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(new_n507_), .Z(new_n550_));
  XNOR2_X1  g349(.A(G127gat), .B(G155gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT16), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(G183gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(G211gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT17), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n550_), .B1(KEYINPUT76), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(KEYINPUT76), .B2(new_n555_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n554_), .A2(KEYINPUT17), .B1(new_n549_), .B2(new_n499_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n549_), .A2(new_n499_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n558_), .B(new_n559_), .C1(KEYINPUT17), .C2(new_n554_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n547_), .A2(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n483_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(G1gat), .B1(new_n564_), .B2(new_n325_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n457_), .A2(new_n482_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n208_), .B1(new_n279_), .B2(new_n269_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT37), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n281_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n281_), .A2(new_n569_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n561_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n524_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n546_), .B(KEYINPUT79), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n566_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(new_n526_), .A3(new_n324_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT104), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT38), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(KEYINPUT104), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n565_), .B1(new_n581_), .B2(new_n582_), .ZN(G1324gat));
  NAND3_X1  g382(.A1(new_n395_), .A2(new_n400_), .A3(new_n403_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n576_), .A2(new_n527_), .A3(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n566_), .A2(new_n282_), .A3(new_n584_), .A4(new_n562_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(G8gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT106), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT106), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n590_), .A3(G8gat), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n588_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n589_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n585_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT40), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(KEYINPUT40), .B(new_n585_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(G1325gat));
  INV_X1    g397(.A(G15gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n563_), .B2(new_n454_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT41), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n576_), .A2(new_n599_), .A3(new_n454_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1326gat));
  INV_X1    g402(.A(G22gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n479_), .B(KEYINPUT107), .Z(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n563_), .B2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT42), .Z(new_n607_));
  NAND3_X1  g406(.A1(new_n576_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1327gat));
  INV_X1    g408(.A(new_n561_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n276_), .A2(new_n280_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n566_), .A2(new_n575_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT109), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT109), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n566_), .A2(new_n615_), .A3(new_n575_), .A4(new_n612_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(G29gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n324_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n547_), .A2(new_n610_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT43), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n569_), .B(new_n611_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n566_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  AOI211_X1 g423(.A(KEYINPUT43), .B(new_n624_), .C1(new_n457_), .C2(new_n482_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n620_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT44), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT44), .B(new_n620_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n324_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT108), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(new_n631_), .A3(G29gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n630_), .B2(G29gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n619_), .B1(new_n632_), .B2(new_n633_), .ZN(G1328gat));
  AOI21_X1  g433(.A(new_n404_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n629_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G36gat), .ZN(new_n637_));
  INV_X1    g436(.A(G36gat), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n614_), .A2(new_n638_), .A3(new_n584_), .A4(new_n616_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT45), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n637_), .A2(KEYINPUT46), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT46), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT45), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n639_), .B(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n638_), .B1(new_n635_), .B2(new_n629_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(new_n646_), .ZN(G1329gat));
  NAND3_X1  g446(.A1(new_n614_), .A2(new_n454_), .A3(new_n616_), .ZN(new_n648_));
  INV_X1    g447(.A(G43gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n628_), .A2(G43gat), .A3(new_n454_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n629_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT47), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT47), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n655_), .B(new_n650_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1330gat));
  AND4_X1   g456(.A1(G50gat), .A2(new_n628_), .A3(new_n479_), .A4(new_n629_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G50gat), .B1(new_n617_), .B2(new_n605_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1331gat));
  AND3_X1   g459(.A1(new_n573_), .A2(new_n610_), .A3(new_n574_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n483_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n325_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n524_), .A2(new_n546_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n566_), .A2(new_n572_), .A3(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(G1332gat));
  INV_X1    g467(.A(G64gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n662_), .B2(new_n584_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT48), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n666_), .A2(new_n669_), .A3(new_n584_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1333gat));
  INV_X1    g472(.A(G71gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n662_), .B2(new_n454_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT49), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n454_), .A2(new_n674_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT110), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n666_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1334gat));
  INV_X1    g479(.A(G78gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n662_), .B2(new_n605_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT50), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n666_), .A2(new_n681_), .A3(new_n605_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1335gat));
  NAND2_X1  g484(.A1(new_n665_), .A2(new_n561_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G85gat), .B1(new_n688_), .B2(new_n325_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n665_), .A2(new_n612_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n566_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n215_), .A3(new_n324_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n689_), .A2(new_n693_), .ZN(G1336gat));
  OAI21_X1  g493(.A(G92gat), .B1(new_n688_), .B2(new_n404_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n692_), .A2(new_n216_), .A3(new_n584_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1337gat));
  OAI21_X1  g496(.A(G99gat), .B1(new_n688_), .B2(new_n481_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n454_), .A2(new_n223_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n691_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g500(.A1(new_n692_), .A2(new_n224_), .A3(new_n479_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n479_), .B(new_n687_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT52), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(G106gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G106gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT53), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT53), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n709_), .B(new_n702_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1339gat));
  INV_X1    g510(.A(KEYINPUT120), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT54), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n522_), .A2(new_n523_), .A3(new_n574_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n572_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n572_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n532_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n544_), .B1(new_n536_), .B2(new_n534_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT115), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n543_), .B2(new_n539_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n519_), .B2(new_n517_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT56), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n518_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n510_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n510_), .A2(KEYINPUT113), .A3(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n510_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n497_), .A2(new_n505_), .A3(new_n500_), .A4(new_n509_), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n739_), .A2(KEYINPUT55), .B1(new_n740_), .B2(new_n502_), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n728_), .B(new_n731_), .C1(new_n738_), .C2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(KEYINPUT55), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n502_), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n498_), .A2(new_n504_), .B1(new_n250_), .B2(new_n508_), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n735_), .B(new_n732_), .C1(new_n745_), .C2(new_n506_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT113), .B1(new_n510_), .B2(new_n733_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n743_), .B(new_n744_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT56), .B1(new_n748_), .B2(new_n516_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT114), .B1(new_n748_), .B2(new_n730_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n742_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n519_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n546_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n727_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT57), .B1(new_n756_), .B2(new_n611_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n748_), .A2(new_n730_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n728_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n748_), .A2(new_n516_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n729_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n731_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT114), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n761_), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n726_), .B1(new_n764_), .B2(new_n754_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n611_), .A2(KEYINPUT57), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n725_), .A2(new_n752_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT58), .B(new_n767_), .C1(new_n749_), .C2(new_n762_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n622_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n518_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n758_), .B1(new_n772_), .B2(KEYINPUT56), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n773_), .B2(new_n767_), .ZN(new_n774_));
  OAI22_X1  g573(.A1(new_n765_), .A2(new_n766_), .B1(new_n769_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n561_), .B1(new_n757_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT119), .ZN(new_n777_));
  INV_X1    g576(.A(new_n766_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n749_), .A2(new_n750_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n755_), .B1(new_n779_), .B2(new_n763_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n780_), .B2(new_n726_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n768_), .A2(new_n622_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n774_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI22_X1  g583(.A1(KEYINPUT114), .A2(new_n762_), .B1(new_n772_), .B2(KEYINPUT56), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n754_), .B1(new_n785_), .B2(new_n742_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n281_), .B1(new_n786_), .B2(new_n727_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n781_), .B(new_n784_), .C1(new_n787_), .C2(KEYINPUT57), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n561_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n720_), .B1(new_n777_), .B2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n440_), .A2(new_n324_), .A3(new_n442_), .A4(new_n454_), .ZN(new_n792_));
  OR3_X1    g591(.A1(new_n792_), .A2(new_n584_), .A3(KEYINPUT117), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT117), .B1(new_n792_), .B2(new_n584_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(KEYINPUT59), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n712_), .B1(new_n791_), .B2(new_n797_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n717_), .A2(new_n719_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n756_), .A2(new_n778_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n765_), .B2(new_n281_), .ZN(new_n802_));
  AOI211_X1 g601(.A(KEYINPUT119), .B(new_n610_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n789_), .B1(new_n788_), .B2(new_n561_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT120), .A3(new_n796_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n610_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n720_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT59), .B1(new_n808_), .B2(new_n795_), .ZN(new_n809_));
  INV_X1    g608(.A(G113gat), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n574_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n798_), .A2(new_n806_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n795_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n546_), .C1(new_n720_), .C2(new_n807_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n814_), .A2(KEYINPUT118), .A3(new_n810_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT118), .B1(new_n814_), .B2(new_n810_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n812_), .A2(KEYINPUT121), .A3(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1340gat));
  NAND3_X1  g621(.A1(new_n798_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n808_), .A2(new_n795_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n524_), .A2(G120gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(KEYINPUT60), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n573_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G120gat), .B1(new_n823_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n561_), .A2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n798_), .A2(new_n806_), .A3(new_n809_), .A4(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n824_), .A2(new_n610_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT122), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT122), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n832_), .A2(new_n837_), .A3(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1342gat));
  OAI21_X1  g638(.A(G134gat), .B1(new_n823_), .B2(new_n624_), .ZN(new_n840_));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n824_), .A2(new_n841_), .A3(new_n283_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1343gat));
  NAND2_X1  g642(.A1(new_n799_), .A2(new_n776_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n404_), .A2(new_n324_), .A3(new_n456_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G141gat), .B1(new_n850_), .B2(new_n753_), .ZN(new_n851_));
  INV_X1    g650(.A(G141gat), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n852_), .B(new_n546_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1344gat));
  OAI21_X1  g653(.A(G148gat), .B1(new_n850_), .B2(new_n524_), .ZN(new_n855_));
  INV_X1    g654(.A(G148gat), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(new_n573_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1345gat));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n850_), .B2(new_n561_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n859_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n610_), .B(new_n861_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1346gat));
  INV_X1    g662(.A(new_n849_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n624_), .B1(new_n864_), .B2(new_n847_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n283_), .A2(new_n205_), .ZN(new_n866_));
  OAI22_X1  g665(.A1(new_n865_), .A2(new_n205_), .B1(new_n850_), .B2(new_n866_), .ZN(G1347gat));
  NOR2_X1   g666(.A1(new_n404_), .A2(new_n324_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n454_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n605_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n805_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT124), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n805_), .A2(new_n873_), .A3(new_n870_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n872_), .A2(new_n337_), .A3(new_n546_), .A4(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G169gat), .B1(new_n871_), .B2(new_n753_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n876_), .A2(KEYINPUT62), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(KEYINPUT62), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n875_), .B1(new_n877_), .B2(new_n878_), .ZN(G1348gat));
  NAND2_X1  g678(.A1(new_n844_), .A2(new_n480_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n880_), .A2(new_n338_), .A3(new_n524_), .A4(new_n869_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n872_), .A2(new_n573_), .A3(new_n874_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n338_), .ZN(G1349gat));
  AND2_X1   g682(.A1(new_n872_), .A2(new_n874_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n561_), .A2(new_n341_), .ZN(new_n885_));
  OR3_X1    g684(.A1(new_n880_), .A2(new_n561_), .A3(new_n869_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n884_), .A2(new_n885_), .B1(new_n326_), .B2(new_n886_), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n872_), .A2(new_n622_), .A3(new_n874_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G190gat), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n872_), .A2(new_n283_), .A3(new_n342_), .A4(new_n874_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1351gat));
  AND2_X1   g690(.A1(new_n868_), .A2(new_n456_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n844_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n546_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g695(.A1(new_n893_), .A2(new_n524_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1353gat));
  AOI21_X1  g698(.A(new_n561_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n894_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT126), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n901_), .A2(new_n902_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n901_), .A2(new_n904_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(G1354gat));
  OR3_X1    g707(.A1(new_n893_), .A2(G218gat), .A3(new_n282_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G218gat), .B1(new_n893_), .B2(new_n624_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1355gat));
endmodule


