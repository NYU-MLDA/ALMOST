//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT22), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT89), .B1(new_n203_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(KEYINPUT22), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT89), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(G176gat), .B1(new_n206_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n214_), .B(new_n215_), .C1(G183gat), .C2(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT90), .B1(new_n211_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n209_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT90), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n219_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n214_), .A2(new_n215_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT87), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT24), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT87), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n227_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n204_), .A2(new_n220_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n217_), .B(new_n235_), .C1(new_n229_), .C2(new_n231_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G183gat), .ZN(new_n239_));
  INV_X1    g038(.A(G183gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT25), .ZN(new_n241_));
  INV_X1    g040(.A(G190gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT26), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT26), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G190gat), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n239_), .A2(new_n241_), .A3(new_n243_), .A4(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n236_), .A2(new_n237_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n237_), .B1(new_n236_), .B2(new_n246_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n234_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n226_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G211gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(G218gat), .ZN(new_n252_));
  INV_X1    g051(.A(G218gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n253_), .A2(G211gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT84), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(G211gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(G218gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261_));
  INV_X1    g060(.A(G197gat), .ZN(new_n262_));
  INV_X1    g061(.A(G204gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G197gat), .A2(G204gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n260_), .A2(new_n261_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n258_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT83), .B1(new_n264_), .B2(new_n265_), .ZN(new_n271_));
  OAI22_X1  g070(.A1(new_n269_), .A2(new_n270_), .B1(new_n271_), .B2(new_n261_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT83), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n266_), .A2(new_n273_), .A3(new_n261_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n272_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(G197gat), .A2(G204gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G197gat), .A2(G204gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n273_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n255_), .A2(new_n259_), .B1(new_n280_), .B2(KEYINPUT21), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT85), .B1(new_n281_), .B2(new_n274_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n268_), .B1(new_n277_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n250_), .A2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n276_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(KEYINPUT85), .A3(new_n274_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n267_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT77), .B1(new_n288_), .B2(G169gat), .ZN(new_n289_));
  AND2_X1   g088(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n290_));
  NOR2_X1   g089(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n291_));
  OAI211_X1 g090(.A(KEYINPUT77), .B(G169gat), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n220_), .B(new_n207_), .C1(new_n289_), .C2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n216_), .A2(KEYINPUT78), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n216_), .A2(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n217_), .A2(KEYINPUT24), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT74), .B1(new_n298_), .B2(new_n233_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n235_), .A2(new_n300_), .A3(KEYINPUT24), .A4(new_n217_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT73), .B1(new_n240_), .B2(KEYINPUT25), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT26), .B(G190gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n303_), .B(new_n304_), .C1(new_n305_), .C2(KEYINPUT73), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT75), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n302_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n227_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n287_), .A2(new_n297_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT19), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n303_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n239_), .A2(new_n241_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n317_), .A2(new_n320_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n311_), .B1(new_n321_), .B2(new_n309_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n310_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n297_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n283_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT20), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n316_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n236_), .A2(new_n246_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT88), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n236_), .A2(new_n237_), .A3(new_n246_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n332_), .A2(new_n234_), .B1(new_n219_), .B2(new_n225_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n328_), .B1(new_n333_), .B2(new_n287_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n314_), .A2(new_n316_), .B1(new_n325_), .B2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G8gat), .B(G36gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n335_), .B(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(KEYINPUT27), .ZN(new_n343_));
  INV_X1    g142(.A(new_n316_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n284_), .A2(new_n313_), .A3(KEYINPUT20), .A4(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n211_), .A2(new_n218_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n332_), .B2(new_n234_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n326_), .B1(new_n347_), .B2(new_n287_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n344_), .B1(new_n348_), .B2(new_n325_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n345_), .B1(new_n349_), .B2(KEYINPUT96), .ZN(new_n350_));
  INV_X1    g149(.A(new_n346_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n249_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT20), .B1(new_n283_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n285_), .A2(new_n286_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n297_), .A2(new_n312_), .B1(new_n354_), .B2(new_n268_), .ZN(new_n355_));
  OAI211_X1 g154(.A(KEYINPUT96), .B(new_n316_), .C1(new_n353_), .C2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n341_), .B1(new_n350_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT97), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT20), .B1(new_n333_), .B2(new_n287_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n324_), .A2(new_n283_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n316_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n334_), .A2(new_n325_), .ZN(new_n364_));
  AND4_X1   g163(.A1(new_n359_), .A2(new_n363_), .A3(new_n340_), .A4(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n358_), .B(KEYINPUT27), .C1(new_n360_), .C2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT98), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n316_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT96), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n356_), .A3(new_n345_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n368_), .B1(new_n372_), .B2(new_n341_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n363_), .A2(new_n340_), .A3(new_n364_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT97), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n335_), .A2(new_n359_), .A3(new_n340_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT98), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n373_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n343_), .B1(new_n367_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n381_));
  INV_X1    g180(.A(G141gat), .ZN(new_n382_));
  INV_X1    g181(.A(G148gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G141gat), .A2(G148gat), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n385_), .A2(KEYINPUT80), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(KEYINPUT80), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n384_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G155gat), .B(G162gat), .Z(new_n389_));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT2), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n385_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n394_), .A2(new_n396_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n389_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n392_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(KEYINPUT29), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT82), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT86), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n402_), .A2(new_n404_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n405_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n388_), .A2(new_n391_), .B1(new_n399_), .B2(new_n389_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n283_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G22gat), .B(G50gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n419_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(G15gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT30), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n324_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G127gat), .B(G134gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G113gat), .B(G120gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(KEYINPUT79), .A3(new_n431_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n427_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438_));
  INV_X1    g237(.A(G43gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT31), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n437_), .B(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G225gat), .A2(G233gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n416_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n416_), .A2(new_n448_), .A3(new_n432_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n435_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT79), .B1(new_n430_), .B2(new_n431_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n401_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n416_), .B2(new_n432_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n444_), .B(new_n447_), .C1(new_n454_), .C2(new_n446_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n416_), .A2(new_n448_), .A3(new_n432_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n453_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n456_), .B1(new_n457_), .B2(new_n445_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n443_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G57gat), .B(G85gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT94), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G1gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n461_), .B(KEYINPUT94), .ZN(new_n465_));
  INV_X1    g264(.A(G1gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n468_));
  INV_X1    g267(.A(G29gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n464_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n460_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n455_), .A2(new_n473_), .A3(new_n459_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n442_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n380_), .A2(new_n422_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n420_), .A2(new_n421_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT95), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484_));
  OR3_X1    g283(.A1(new_n476_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n476_), .B2(new_n484_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n443_), .B(new_n447_), .C1(new_n454_), .C2(new_n446_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n473_), .B1(new_n458_), .B2(new_n444_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n476_), .B1(new_n489_), .B2(new_n484_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n342_), .A2(new_n485_), .A3(new_n486_), .A4(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n340_), .A2(KEYINPUT32), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n335_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n372_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n477_), .B(new_n493_), .C1(new_n494_), .C2(new_n492_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n482_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n422_), .A2(new_n477_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n380_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n481_), .B1(new_n498_), .B2(new_n442_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT6), .ZN(new_n502_));
  INV_X1    g301(.A(G99gat), .ZN(new_n503_));
  INV_X1    g302(.A(G106gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n504_), .A3(KEYINPUT64), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT7), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n507_), .A2(new_n503_), .A3(new_n504_), .A4(KEYINPUT64), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n502_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G85gat), .B(G92gat), .Z(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT65), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT8), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(KEYINPUT65), .A3(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n504_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT9), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(G85gat), .A3(G92gat), .ZN(new_n520_));
  AND4_X1   g319(.A1(new_n502_), .A2(new_n517_), .A3(new_n518_), .A4(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n526_));
  XOR2_X1   g325(.A(G71gat), .B(G78gat), .Z(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n526_), .A2(new_n527_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n500_), .B1(new_n523_), .B2(new_n531_), .ZN(new_n532_));
  AOI211_X1 g331(.A(KEYINPUT12), .B(new_n530_), .C1(new_n515_), .C2(new_n522_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n515_), .A2(new_n530_), .A3(new_n522_), .ZN(new_n535_));
  INV_X1    g334(.A(G230gat), .ZN(new_n536_));
  INV_X1    g335(.A(G233gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT66), .B1(new_n534_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n523_), .A2(new_n531_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n535_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n538_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n540_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n545_), .B(new_n546_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n541_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G120gat), .B(G148gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT5), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n552_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n541_), .A2(new_n544_), .A3(new_n547_), .A4(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n553_), .A2(KEYINPUT13), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT13), .B1(new_n553_), .B2(new_n555_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G29gat), .B(G36gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G43gat), .B(G50gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT15), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G15gat), .B(G22gat), .ZN(new_n564_));
  INV_X1    g363(.A(G8gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT14), .B1(new_n466_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G1gat), .B(G8gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  OR2_X1    g368(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n561_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n572_), .B(KEYINPUT71), .Z(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(KEYINPUT70), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n569_), .A2(new_n561_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n574_), .B1(new_n577_), .B2(new_n572_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G113gat), .B(G141gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT72), .ZN(new_n580_));
  XOR2_X1   g379(.A(G169gat), .B(G197gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n578_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n558_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n515_), .A2(new_n522_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n561_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n563_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n523_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n563_), .B1(new_n515_), .B2(new_n522_), .ZN(new_n595_));
  OAI211_X1 g394(.A(KEYINPUT35), .B(new_n594_), .C1(new_n595_), .C2(KEYINPUT68), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n590_), .A2(new_n596_), .B1(KEYINPUT36), .B2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n595_), .B1(new_n561_), .B2(new_n586_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n594_), .A2(KEYINPUT35), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT68), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n589_), .B2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n594_), .A2(KEYINPUT35), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n600_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n599_), .A2(KEYINPUT36), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n608_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n600_), .A2(new_n606_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(KEYINPUT69), .A2(KEYINPUT37), .ZN(new_n613_));
  OR2_X1    g412(.A1(KEYINPUT69), .A2(KEYINPUT37), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n609_), .A2(KEYINPUT69), .A3(KEYINPUT37), .A4(new_n611_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n569_), .B(new_n530_), .Z(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  XOR2_X1   g420(.A(G127gat), .B(G155gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT16), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n620_), .A2(new_n621_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(KEYINPUT17), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n620_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n617_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n499_), .A2(new_n585_), .A3(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT99), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(KEYINPUT99), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n634_), .A2(new_n466_), .A3(new_n477_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n636_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(KEYINPUT38), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n584_), .A2(KEYINPUT101), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n558_), .A2(new_n641_), .A3(new_n583_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n612_), .B(KEYINPUT102), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n499_), .A2(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n643_), .A2(new_n646_), .A3(new_n629_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n478_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n639_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT38), .B1(new_n637_), .B2(new_n638_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1324gat));
  INV_X1    g451(.A(new_n380_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n634_), .A2(new_n565_), .A3(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT103), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n565_), .B1(new_n647_), .B2(new_n653_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT39), .Z(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(G1325gat));
  AOI21_X1  g459(.A(new_n424_), .B1(new_n647_), .B2(new_n442_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT41), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n634_), .A2(new_n424_), .A3(new_n442_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n647_), .B2(new_n482_), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n634_), .A2(new_n665_), .A3(new_n482_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(new_n629_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n645_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n499_), .A2(new_n672_), .A3(new_n585_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n477_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n671_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n499_), .B2(new_n617_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n342_), .A2(KEYINPUT27), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n373_), .A2(new_n378_), .A3(new_n377_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n378_), .B1(new_n373_), .B2(new_n377_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n497_), .B(new_n679_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n363_), .A2(new_n364_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n341_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n490_), .A2(new_n486_), .A3(new_n374_), .A4(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n485_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n495_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n422_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n442_), .B1(new_n682_), .B2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n422_), .B(new_n679_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n479_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n677_), .B(new_n617_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n676_), .B1(new_n678_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n676_), .C1(new_n678_), .C2(new_n693_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n478_), .A2(new_n469_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n675_), .B1(new_n698_), .B2(new_n699_), .ZN(G1328gat));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n380_), .B(KEYINPUT106), .Z(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT108), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n674_), .A2(new_n701_), .A3(new_n702_), .A4(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n704_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n702_), .A2(new_n701_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n673_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n696_), .A2(new_n653_), .A3(new_n697_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G36gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT110), .B1(new_n711_), .B2(KEYINPUT109), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT111), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  INV_X1    g513(.A(new_n711_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT110), .B(new_n718_), .C1(new_n711_), .C2(KEYINPUT109), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n713_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n717_), .B1(new_n713_), .B2(new_n719_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  NAND3_X1  g521(.A1(new_n698_), .A2(G43gat), .A3(new_n442_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n442_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n439_), .B1(new_n673_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n674_), .B2(new_n482_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n482_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n698_), .B2(new_n730_), .ZN(G1331gat));
  NOR2_X1   g530(.A1(new_n558_), .A2(new_n583_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n499_), .A2(new_n671_), .A3(new_n645_), .A4(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT113), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n478_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n499_), .A2(new_n732_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n630_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n477_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n743_), .A3(new_n702_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n734_), .A2(new_n702_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G64gat), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT48), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(KEYINPUT48), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1333gat));
  OR3_X1    g548(.A1(new_n738_), .A2(G71gat), .A3(new_n724_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G71gat), .B1(new_n735_), .B2(new_n724_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT49), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(KEYINPUT49), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1334gat));
  OR3_X1    g553(.A1(new_n738_), .A2(G78gat), .A3(new_n422_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G78gat), .B1(new_n735_), .B2(new_n422_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(KEYINPUT50), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT50), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n755_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  INV_X1    g558(.A(G85gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n737_), .A2(new_n672_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n478_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT114), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n629_), .B(new_n732_), .C1(new_n678_), .C2(new_n693_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT115), .Z(new_n765_));
  NOR2_X1   g564(.A1(new_n478_), .A2(new_n760_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT116), .ZN(G1336gat));
  INV_X1    g567(.A(new_n761_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G92gat), .B1(new_n769_), .B2(new_n653_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n702_), .A2(G92gat), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT117), .Z(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n765_), .B2(new_n772_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT118), .Z(G1337gat));
  AND3_X1   g573(.A1(new_n769_), .A2(new_n516_), .A3(new_n442_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n765_), .A2(new_n442_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(G99gat), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n504_), .A3(new_n482_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n764_), .A2(new_n422_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G106gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g584(.A1(new_n690_), .A2(new_n478_), .A3(new_n724_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n615_), .A2(new_n616_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n578_), .A2(new_n582_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n573_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n570_), .A2(new_n571_), .A3(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n582_), .B(new_n791_), .C1(new_n577_), .C2(new_n790_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n555_), .A2(new_n789_), .A3(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n534_), .A2(new_n540_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n535_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n794_), .A2(KEYINPUT55), .B1(new_n795_), .B2(new_n538_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n541_), .A2(new_n547_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(KEYINPUT55), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n552_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n793_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n788_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n793_), .B(KEYINPUT58), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n798_), .A2(new_n552_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n811_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n793_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n803_), .A2(new_n806_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n583_), .A2(new_n555_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n789_), .A2(new_n792_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n645_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n813_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n818_), .A2(new_n819_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n629_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n583_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n671_), .A2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT119), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(new_n788_), .A3(new_n558_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT54), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n787_), .B1(new_n823_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829_), .B2(new_n583_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n813_), .A2(new_n820_), .A3(KEYINPUT121), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT121), .B1(new_n813_), .B2(new_n820_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n822_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT122), .B1(new_n835_), .B2(new_n671_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n822_), .B1(new_n821_), .B2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n813_), .A2(new_n820_), .A3(KEYINPUT121), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n671_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n836_), .A2(new_n842_), .A3(new_n828_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n787_), .A2(KEYINPUT59), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n832_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n824_), .A2(KEYINPUT123), .ZN(new_n846_));
  MUX2_X1   g645(.A(KEYINPUT123), .B(new_n846_), .S(G113gat), .Z(new_n847_));
  AOI21_X1  g646(.A(new_n830_), .B1(new_n845_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n558_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n829_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n849_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n558_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n855_));
  OAI21_X1  g654(.A(G120gat), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT124), .B(new_n853_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n851_), .B1(new_n856_), .B2(new_n857_), .ZN(G1341gat));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n829_), .A2(new_n859_), .A3(new_n671_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n845_), .A2(new_n671_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n859_), .ZN(G1342gat));
  INV_X1    g661(.A(G134gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n829_), .A2(new_n863_), .A3(new_n644_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n845_), .A2(new_n617_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1343gat));
  AOI21_X1  g665(.A(new_n442_), .B1(new_n823_), .B2(new_n828_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n702_), .A2(new_n478_), .A3(new_n422_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n824_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n382_), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n558_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n383_), .ZN(G1345gat));
  NOR2_X1   g672(.A1(new_n869_), .A2(new_n629_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  OAI21_X1  g675(.A(G162gat), .B1(new_n869_), .B2(new_n788_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n645_), .A2(G162gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n869_), .B2(new_n878_), .ZN(G1347gat));
  NAND2_X1  g678(.A1(new_n702_), .A2(new_n480_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT125), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n482_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n828_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n835_), .A2(KEYINPUT122), .A3(new_n671_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n583_), .B(new_n882_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n885_), .A2(new_n886_), .A3(G169gat), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n843_), .A2(new_n882_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n888_), .B(new_n583_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n886_), .B1(new_n885_), .B2(G169gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(G1348gat));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n852_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n482_), .B1(new_n823_), .B2(new_n828_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n881_), .A2(new_n220_), .A3(new_n558_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n892_), .A2(new_n220_), .B1(new_n893_), .B2(new_n894_), .ZN(G1349gat));
  NOR2_X1   g694(.A1(new_n881_), .A2(new_n629_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G183gat), .B1(new_n893_), .B2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n629_), .A2(new_n305_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n888_), .B2(new_n898_), .ZN(G1350gat));
  NAND2_X1  g698(.A1(new_n888_), .A2(new_n617_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(G190gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n888_), .A2(new_n304_), .A3(new_n644_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1351gat));
  AND2_X1   g702(.A1(new_n702_), .A2(new_n497_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n867_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n824_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n262_), .ZN(G1352gat));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n558_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n263_), .ZN(G1353gat));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n671_), .B1(new_n910_), .B2(new_n251_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT126), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n867_), .A2(new_n904_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n251_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1354gat));
  OAI21_X1  g714(.A(G218gat), .B1(new_n905_), .B2(new_n788_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n644_), .A2(new_n253_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n905_), .B2(new_n917_), .ZN(G1355gat));
endmodule


