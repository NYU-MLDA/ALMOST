//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT86), .B(G197gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G211gat), .B(G218gat), .Z(new_n210_));
  NAND2_X1  g009(.A1(new_n203_), .A2(new_n205_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n208_), .B1(G197gat), .B2(G204gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(KEYINPUT21), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n207_), .A2(KEYINPUT87), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n204_), .A2(new_n206_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT29), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT3), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT2), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(KEYINPUT1), .B2(new_n228_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(KEYINPUT1), .B2(new_n228_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n223_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n225_), .A3(new_n234_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  OAI22_X1  g035(.A1(new_n215_), .A2(new_n221_), .B1(new_n222_), .B2(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(G228gat), .A2(G233gat), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n241_), .A2(KEYINPUT88), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(KEYINPUT88), .ZN(new_n243_));
  OAI211_X1 g042(.A(KEYINPUT89), .B(new_n202_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(new_n222_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G22gat), .B(G50gat), .Z(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n241_), .A2(new_n202_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT90), .ZN(new_n252_));
  OR3_X1    g051(.A1(new_n241_), .A2(KEYINPUT90), .A3(new_n202_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n244_), .A2(new_n249_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n242_), .A2(new_n243_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT89), .B1(new_n255_), .B2(new_n202_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n241_), .A2(new_n202_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n251_), .A2(new_n257_), .ZN(new_n258_));
  OAI22_X1  g057(.A1(new_n254_), .A2(new_n256_), .B1(new_n258_), .B2(new_n249_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n217_), .A2(new_n220_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n216_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n214_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT82), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n266_), .A2(KEYINPUT24), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(KEYINPUT24), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT23), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT25), .B(G183gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n267_), .A2(new_n269_), .A3(new_n271_), .A4(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n271_), .B1(G183gat), .B2(G190gat), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  INV_X1    g076(.A(G169gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT83), .B1(new_n278_), .B2(KEYINPUT22), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT22), .B(G169gat), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n277_), .B(new_n279_), .C1(new_n280_), .C2(KEYINPUT83), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n276_), .A2(new_n281_), .A3(new_n268_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n260_), .B1(new_n264_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT93), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G226gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n265_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n271_), .B1(KEYINPUT24), .B2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n291_), .A2(KEYINPUT92), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(KEYINPUT92), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n292_), .A2(new_n274_), .A3(new_n269_), .A4(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n280_), .A2(new_n277_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n276_), .A2(new_n268_), .A3(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n263_), .A2(new_n214_), .A3(new_n294_), .A4(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n284_), .A2(new_n285_), .A3(new_n289_), .A4(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n283_), .B1(new_n215_), .B2(new_n221_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n297_), .A2(new_n299_), .A3(KEYINPUT20), .A4(new_n289_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT93), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n294_), .A2(new_n296_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n260_), .B1(new_n264_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n283_), .B2(new_n264_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n288_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G8gat), .B(G36gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(G64gat), .B(G92gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n302_), .A2(new_n306_), .A3(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n305_), .A2(new_n289_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n284_), .A2(new_n288_), .A3(new_n297_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n313_), .A3(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(KEYINPUT27), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n259_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n283_), .B(KEYINPUT30), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G71gat), .B(G99gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(G43gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G227gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(G15gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n328_), .B(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n326_), .B(new_n332_), .Z(new_n333_));
  AND2_X1   g132(.A1(new_n333_), .A2(KEYINPUT84), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(KEYINPUT84), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G127gat), .B(G134gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G113gat), .B(G120gat), .Z(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n336_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT31), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n334_), .A2(new_n335_), .A3(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n333_), .A2(KEYINPUT84), .A3(new_n343_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n342_), .A2(KEYINPUT95), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n342_), .A2(KEYINPUT95), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n236_), .B(KEYINPUT96), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n339_), .A2(new_n341_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT95), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n231_), .A2(new_n235_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT96), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n353_), .B2(new_n351_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n350_), .B(KEYINPUT4), .C1(new_n354_), .C2(new_n356_), .ZN(new_n357_));
  OR3_X1    g156(.A1(new_n236_), .A2(KEYINPUT4), .A3(new_n342_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n347_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT0), .ZN(new_n362_));
  INV_X1    g161(.A(G57gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(G85gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n347_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n356_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n353_), .B2(new_n352_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n369_), .B2(new_n350_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n360_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n366_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n359_), .B2(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n346_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n325_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT101), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n312_), .A2(KEYINPUT32), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n302_), .A2(new_n306_), .A3(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n319_), .A2(KEYINPUT32), .A3(new_n312_), .A4(new_n320_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n375_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT100), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT97), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  OR3_X1    g186(.A1(new_n374_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n374_), .B2(new_n387_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n367_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n347_), .B1(new_n369_), .B2(new_n350_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n366_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT98), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT98), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n395_), .B(new_n366_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n374_), .A2(new_n387_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n397_), .A2(new_n314_), .A3(new_n315_), .A4(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT99), .B1(new_n390_), .B2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n314_), .A2(new_n315_), .A3(new_n398_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT99), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n388_), .A2(new_n389_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .A4(new_n397_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n385_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n379_), .B1(new_n405_), .B2(new_n259_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n400_), .A2(new_n404_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n385_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n259_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(KEYINPUT101), .A3(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n323_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n375_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n378_), .B1(new_n415_), .B2(new_n346_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G1gat), .B(G8gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n418_), .B(KEYINPUT78), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G1gat), .ZN(new_n421_));
  INV_X1    g220(.A(G8gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT14), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G22gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G15gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n330_), .A2(G22gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT77), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(KEYINPUT77), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n420_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n419_), .A2(new_n429_), .A3(new_n428_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G29gat), .B(G36gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G43gat), .B(G50gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n417_), .B1(new_n433_), .B2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT79), .A4(new_n436_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n433_), .A2(new_n437_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G229gat), .A2(G233gat), .ZN(new_n443_));
  OR3_X1    g242(.A1(new_n442_), .A2(KEYINPUT80), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT80), .B1(new_n442_), .B2(new_n443_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n436_), .B(KEYINPUT15), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n433_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n440_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n443_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n444_), .A2(new_n445_), .A3(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G113gat), .B(G141gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT81), .ZN(new_n453_));
  XOR2_X1   g252(.A(G169gat), .B(G197gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n455_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n444_), .A2(new_n445_), .A3(new_n450_), .A4(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G230gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT64), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT65), .ZN(new_n463_));
  AND2_X1   g262(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G106gat), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n463_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NOR4_X1   g267(.A1(new_n464_), .A2(new_n465_), .A3(KEYINPUT65), .A4(G106gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT68), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT68), .ZN(new_n477_));
  NAND3_X1  g276(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n473_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G85gat), .A2(G92gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G85gat), .A2(G92gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT66), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n483_), .B2(KEYINPUT9), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT9), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(KEYINPUT66), .A3(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n484_), .A2(KEYINPUT67), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT67), .B1(new_n484_), .B2(new_n486_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n470_), .B(new_n480_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT7), .ZN(new_n490_));
  INV_X1    g289(.A(G99gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n467_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n492_), .A2(new_n476_), .A3(new_n478_), .A4(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G85gat), .B(G92gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT69), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(new_n498_), .A3(new_n495_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(KEYINPUT8), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n493_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(new_n473_), .A3(new_n479_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n495_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT8), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n489_), .A2(new_n500_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G71gat), .B(G78gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G57gat), .B(G64gat), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(KEYINPUT11), .B2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n514_));
  INV_X1    g313(.A(new_n509_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n508_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT71), .ZN(new_n519_));
  AND4_X1   g318(.A1(new_n489_), .A2(new_n500_), .A3(new_n516_), .A4(new_n507_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n462_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT72), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT8), .B1(new_n504_), .B2(new_n495_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n499_), .A2(KEYINPUT8), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n526_), .B2(new_n497_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n516_), .B1(new_n527_), .B2(new_n489_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT73), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT12), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n520_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n529_), .A2(KEYINPUT12), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n530_), .B1(new_n518_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n462_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n523_), .A2(KEYINPUT72), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n524_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT5), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G176gat), .B(G204gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n538_), .B(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT13), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT13), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n416_), .A2(new_n460_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT34), .Z(new_n552_));
  NAND2_X1  g351(.A1(new_n508_), .A2(new_n446_), .ZN(new_n553_));
  AOI211_X1 g352(.A(new_n550_), .B(new_n552_), .C1(new_n553_), .C2(KEYINPUT75), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n550_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT74), .Z(new_n556_));
  OAI211_X1 g355(.A(new_n553_), .B(new_n556_), .C1(new_n508_), .C2(new_n437_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n554_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G190gat), .B(G218gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT76), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n558_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n558_), .A2(new_n564_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT37), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n433_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(new_n517_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n576_), .A2(new_n577_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n572_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n578_), .B2(new_n572_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n569_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n549_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n421_), .A3(new_n375_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT38), .ZN(new_n586_));
  INV_X1    g385(.A(new_n568_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n416_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n548_), .A2(new_n460_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n581_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G1gat), .B1(new_n590_), .B2(new_n413_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(G1324gat));
  INV_X1    g391(.A(new_n323_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G8gat), .B1(new_n590_), .B2(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT39), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(KEYINPUT39), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n593_), .A2(G8gat), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n595_), .A2(new_n596_), .B1(new_n584_), .B2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(G1325gat));
  INV_X1    g399(.A(new_n590_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n346_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n330_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT41), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n604_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n584_), .A2(new_n330_), .A3(new_n602_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .ZN(G1326gat));
  OAI21_X1  g407(.A(G22gat), .B1(new_n590_), .B2(new_n410_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT42), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n584_), .A2(new_n424_), .A3(new_n259_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1327gat));
  INV_X1    g411(.A(new_n581_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n549_), .A2(new_n587_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(G29gat), .B1(new_n614_), .B2(new_n375_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT44), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT104), .B1(new_n616_), .B2(KEYINPUT105), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n415_), .A2(new_n346_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n378_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT43), .ZN(new_n621_));
  INV_X1    g420(.A(new_n569_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT43), .B1(new_n416_), .B2(new_n569_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n589_), .A2(new_n613_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n617_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT105), .B1(new_n628_), .B2(KEYINPUT104), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n627_), .B1(new_n629_), .B2(KEYINPUT44), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n375_), .A2(G29gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n615_), .B1(new_n630_), .B2(new_n631_), .ZN(G1328gat));
  INV_X1    g431(.A(KEYINPUT46), .ZN(new_n633_));
  INV_X1    g432(.A(G36gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n630_), .B2(new_n323_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n614_), .A2(new_n634_), .A3(new_n323_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT45), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n633_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n636_), .B(KEYINPUT45), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  AOI211_X1 g440(.A(new_n641_), .B(new_n626_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n616_), .B1(new_n642_), .B2(KEYINPUT105), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n593_), .B1(new_n643_), .B2(new_n627_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n640_), .B(KEYINPUT46), .C1(new_n644_), .C2(new_n634_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(new_n645_), .ZN(G1329gat));
  INV_X1    g445(.A(KEYINPUT47), .ZN(new_n647_));
  INV_X1    g446(.A(G43gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n630_), .B2(new_n602_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n614_), .A2(new_n648_), .A3(new_n602_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n647_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n346_), .B1(new_n643_), .B2(new_n627_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT47), .B(new_n650_), .C1(new_n653_), .C2(new_n648_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1330gat));
  AOI21_X1  g454(.A(G50gat), .B1(new_n614_), .B2(new_n259_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n259_), .A2(G50gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n630_), .B2(new_n657_), .ZN(G1331gat));
  NAND2_X1  g457(.A1(new_n548_), .A2(new_n583_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n460_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n416_), .B(new_n661_), .C1(new_n660_), .C2(new_n659_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n363_), .A3(new_n375_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n548_), .A2(new_n460_), .ZN(new_n664_));
  NOR4_X1   g463(.A1(new_n416_), .A2(new_n587_), .A3(new_n613_), .A4(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(new_n375_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n666_), .B2(new_n363_), .ZN(G1332gat));
  INV_X1    g466(.A(G64gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n665_), .B2(new_n323_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT48), .Z(new_n670_));
  NAND3_X1  g469(.A1(new_n662_), .A2(new_n668_), .A3(new_n323_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1333gat));
  INV_X1    g471(.A(G71gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n662_), .A2(new_n673_), .A3(new_n602_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n665_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G71gat), .B1(new_n675_), .B2(new_n346_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT49), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT49), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(G1334gat));
  INV_X1    g480(.A(G78gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n665_), .B2(new_n259_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT50), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n662_), .A2(new_n682_), .A3(new_n259_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1335gat));
  NAND2_X1  g485(.A1(new_n625_), .A2(KEYINPUT109), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n623_), .A2(new_n624_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n664_), .A2(new_n581_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n687_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n365_), .A3(new_n413_), .ZN(new_n693_));
  NOR4_X1   g492(.A1(new_n416_), .A2(new_n568_), .A3(new_n581_), .A4(new_n664_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G85gat), .B1(new_n694_), .B2(new_n375_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT108), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1336gat));
  OAI21_X1  g496(.A(G92gat), .B1(new_n692_), .B2(new_n593_), .ZN(new_n698_));
  INV_X1    g497(.A(G92gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n694_), .A2(new_n699_), .A3(new_n323_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1337gat));
  OAI21_X1  g500(.A(G99gat), .B1(new_n692_), .B2(new_n346_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n694_), .A2(new_n466_), .A3(new_n602_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT51), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n702_), .A2(new_n706_), .A3(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1338gat));
  NAND2_X1  g507(.A1(new_n691_), .A2(new_n259_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G106gat), .B1(new_n625_), .B2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n711_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n694_), .A2(new_n467_), .A3(new_n259_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n712_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT53), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n712_), .A2(new_n717_), .A3(new_n713_), .A4(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1339gat));
  NAND3_X1  g518(.A1(new_n547_), .A2(new_n583_), .A3(new_n460_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT54), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n533_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n531_), .B1(new_n528_), .B2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n508_), .A2(new_n517_), .A3(new_n531_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n527_), .A2(new_n489_), .A3(new_n516_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n724_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT112), .B1(new_n532_), .B2(new_n534_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n462_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI211_X1 g532(.A(KEYINPUT113), .B(new_n462_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n536_), .A2(KEYINPUT111), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT55), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT55), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n536_), .A2(KEYINPUT111), .A3(new_n737_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n733_), .A2(new_n734_), .A3(new_n736_), .A4(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(KEYINPUT56), .A3(new_n542_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT116), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n739_), .A2(new_n742_), .A3(KEYINPUT56), .A4(new_n542_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n734_), .A2(new_n736_), .A3(new_n738_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n728_), .B1(new_n724_), .B2(new_n727_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n532_), .A2(new_n534_), .A3(KEYINPUT112), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT113), .B1(new_n748_), .B2(new_n462_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n542_), .B1(new_n745_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n744_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT58), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n538_), .A2(new_n543_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n443_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n457_), .B1(new_n449_), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n756_), .B2(new_n442_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n458_), .A2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .A4(new_n759_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n741_), .A2(new_n743_), .B1(new_n751_), .B2(new_n750_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n755_), .A2(new_n759_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT58), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n569_), .B1(new_n760_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT117), .ZN(new_n765_));
  INV_X1    g564(.A(new_n740_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n752_), .A2(KEYINPUT114), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n750_), .A2(new_n768_), .A3(new_n751_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n766_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n459_), .A2(new_n755_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT115), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT114), .B(KEYINPUT56), .C1(new_n739_), .C2(new_n542_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n768_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n740_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n771_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n544_), .A2(new_n759_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n772_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n568_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT57), .A3(new_n568_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n765_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n722_), .B1(new_n786_), .B2(new_n613_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n325_), .A2(new_n413_), .A3(new_n346_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n459_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  INV_X1    g591(.A(G113gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n787_), .A2(new_n460_), .A3(new_n789_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT118), .B1(new_n795_), .B2(G113gat), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n764_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n784_), .A2(new_n798_), .A3(new_n785_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n722_), .B1(new_n799_), .B2(new_n613_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n800_), .A2(KEYINPUT59), .A3(new_n789_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT59), .B1(new_n787_), .B2(new_n789_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT119), .B(KEYINPUT59), .C1(new_n787_), .C2(new_n789_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT120), .B(G113gat), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n460_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n797_), .B1(new_n806_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g608(.A(KEYINPUT60), .ZN(new_n810_));
  INV_X1    g609(.A(G120gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n548_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n790_), .A2(new_n813_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n547_), .B(new_n801_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n811_), .ZN(G1341gat));
  INV_X1    g615(.A(G127gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n790_), .A2(new_n817_), .A3(new_n581_), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n613_), .B(new_n801_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n817_), .ZN(G1342gat));
  INV_X1    g619(.A(G134gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n790_), .A2(new_n821_), .A3(new_n587_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n569_), .B(new_n801_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n821_), .ZN(G1343gat));
  NAND2_X1  g623(.A1(new_n786_), .A2(new_n613_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n722_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NOR4_X1   g626(.A1(new_n410_), .A2(new_n413_), .A3(new_n602_), .A4(new_n323_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n459_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n548_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g633(.A1(new_n829_), .A2(new_n613_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT61), .B(G155gat), .Z(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1346gat));
  OR3_X1    g636(.A1(new_n829_), .A2(G162gat), .A3(new_n568_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G162gat), .B1(new_n829_), .B2(new_n569_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1347gat));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n377_), .A2(new_n259_), .A3(new_n593_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n775_), .A2(new_n776_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n779_), .B1(new_n844_), .B2(KEYINPUT115), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n587_), .B1(new_n845_), .B2(new_n778_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n798_), .B1(new_n846_), .B2(KEYINPUT57), .ZN(new_n847_));
  INV_X1    g646(.A(new_n785_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n613_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n843_), .B1(new_n849_), .B2(new_n826_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n841_), .B1(new_n850_), .B2(new_n459_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n800_), .A2(KEYINPUT121), .A3(new_n460_), .A4(new_n843_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G169gat), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(KEYINPUT123), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n764_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n581_), .B1(new_n858_), .B2(new_n785_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n459_), .B(new_n842_), .C1(new_n859_), .C2(new_n722_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT121), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n849_), .A2(new_n826_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n862_), .A2(new_n841_), .A3(new_n459_), .A4(new_n842_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n278_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n857_), .B1(new_n864_), .B2(new_n854_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n854_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n856_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n850_), .A2(new_n280_), .A3(new_n459_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1348gat));
  AOI21_X1  g668(.A(G176gat), .B1(new_n850_), .B2(new_n548_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n827_), .A2(G176gat), .A3(new_n548_), .A4(new_n842_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(KEYINPUT124), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(KEYINPUT124), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n870_), .B1(new_n872_), .B2(new_n873_), .ZN(G1349gat));
  INV_X1    g673(.A(new_n850_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n875_), .A2(new_n272_), .A3(new_n613_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n787_), .A2(new_n613_), .A3(new_n843_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G183gat), .B1(new_n877_), .B2(new_n878_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n876_), .B1(new_n879_), .B2(new_n880_), .ZN(G1350gat));
  OAI21_X1  g680(.A(G190gat), .B1(new_n875_), .B2(new_n569_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n850_), .A2(new_n587_), .A3(new_n273_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1351gat));
  NOR4_X1   g683(.A1(new_n410_), .A2(new_n593_), .A3(new_n602_), .A4(new_n375_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n827_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n459_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g687(.A(new_n547_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n891_));
  XOR2_X1   g690(.A(new_n890_), .B(new_n891_), .Z(G1353gat));
  NAND2_X1  g691(.A1(new_n827_), .A2(new_n885_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n613_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  AND2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n894_), .B2(new_n895_), .ZN(G1354gat));
  AND3_X1   g697(.A1(new_n886_), .A2(G218gat), .A3(new_n622_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n893_), .A2(KEYINPUT127), .A3(new_n568_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(G218gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT127), .B1(new_n893_), .B2(new_n568_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n901_), .B2(new_n902_), .ZN(G1355gat));
endmodule


