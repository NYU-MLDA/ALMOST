//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT0), .ZN(new_n203_));
  INV_X1    g002(.A(G57gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT102), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G155gat), .B(G162gat), .Z(new_n211_));
  INV_X1    g010(.A(G141gat), .ZN(new_n212_));
  INV_X1    g011(.A(G148gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT93), .ZN(new_n215_));
  AOI22_X1  g014(.A1(KEYINPUT2), .A2(new_n214_), .B1(new_n215_), .B2(KEYINPUT3), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(KEYINPUT3), .B2(new_n215_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n218_), .B(KEYINPUT94), .Z(new_n219_));
  OAI21_X1  g018(.A(new_n211_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n211_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n214_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n212_), .A2(new_n213_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n229_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT101), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT92), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(new_n231_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n227_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT4), .B1(new_n234_), .B2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(KEYINPUT4), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n210_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n227_), .A2(new_n233_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n237_), .B2(new_n227_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(new_n209_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n207_), .B1(new_n241_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n207_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n238_), .A2(KEYINPUT4), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(KEYINPUT4), .B2(new_n243_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n246_), .B(new_n247_), .C1(new_n249_), .C2(new_n210_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G64gat), .B(G92gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n254_), .B(new_n255_), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT32), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT19), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G190gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT86), .B1(new_n263_), .B2(KEYINPUT26), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT25), .B(G183gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G190gat), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n264_), .B(new_n265_), .C1(new_n266_), .C2(KEYINPUT86), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT87), .ZN(new_n268_));
  INV_X1    g067(.A(G183gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT23), .B1(new_n269_), .B2(new_n263_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(G183gat), .A3(G190gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT24), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276_));
  MUX2_X1   g075(.A(new_n275_), .B(KEYINPUT24), .S(new_n276_), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n268_), .A2(new_n273_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n274_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT22), .B(G169gat), .ZN(new_n280_));
  INV_X1    g079(.A(G176gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n272_), .A2(KEYINPUT88), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n270_), .A2(new_n272_), .A3(KEYINPUT88), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n278_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT89), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n278_), .A2(KEYINPUT89), .A3(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G204gat), .ZN(new_n293_));
  OR3_X1    g092(.A1(new_n293_), .A2(KEYINPUT97), .A3(G197gat), .ZN(new_n294_));
  INV_X1    g093(.A(G197gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G204gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT97), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(G197gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT21), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n298_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n300_), .B(new_n301_), .C1(KEYINPUT21), .C2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT98), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n301_), .B(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(KEYINPUT21), .A3(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n292_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT20), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n303_), .A2(new_n306_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n266_), .A2(new_n265_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n277_), .A2(new_n283_), .A3(new_n284_), .A4(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n273_), .B1(G183gat), .B2(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n282_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n309_), .B1(new_n310_), .B2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n262_), .B1(new_n308_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n290_), .A2(new_n291_), .A3(new_n310_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n312_), .A2(KEYINPUT99), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(KEYINPUT99), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n314_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n309_), .B1(new_n321_), .B2(new_n307_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n318_), .A2(new_n262_), .A3(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n259_), .B1(new_n317_), .B2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n262_), .B1(new_n318_), .B2(new_n322_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n310_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n327_));
  OAI211_X1 g126(.A(KEYINPUT20), .B(new_n262_), .C1(new_n321_), .C2(new_n307_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(new_n329_), .A3(new_n258_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n251_), .A2(new_n324_), .A3(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n326_), .A2(new_n329_), .A3(new_n257_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n327_), .A2(new_n328_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n256_), .B1(new_n325_), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n207_), .B1(new_n243_), .B2(new_n210_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT103), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n209_), .B2(new_n249_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n335_), .A2(new_n336_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n332_), .B(new_n334_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT33), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n250_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n241_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n343_), .A2(KEYINPUT33), .A3(new_n246_), .A4(new_n247_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n331_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT96), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n347_), .B(new_n307_), .C1(new_n227_), .C2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G228gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n310_), .A2(KEYINPUT96), .ZN(new_n354_));
  INV_X1    g153(.A(new_n352_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n354_), .B(new_n355_), .C1(new_n348_), .C2(new_n227_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n227_), .A2(new_n348_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G22gat), .B(G50gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(new_n227_), .B2(new_n348_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n362_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n227_), .A2(new_n348_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n358_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n367_), .B2(new_n360_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n357_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n362_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n365_), .A3(new_n360_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n353_), .A4(new_n356_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n346_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT27), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n257_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n325_), .A2(new_n333_), .A3(new_n256_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n373_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n256_), .B1(new_n317_), .B2(new_n323_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(KEYINPUT27), .A3(new_n332_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT104), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n379_), .A2(new_n380_), .A3(new_n382_), .A4(KEYINPUT104), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n375_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G15gat), .B(G43gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n290_), .A2(KEYINPUT30), .A3(new_n291_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT30), .B1(new_n290_), .B2(new_n291_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n391_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n392_), .A3(new_n390_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n389_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n237_), .B(KEYINPUT31), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT91), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n402_), .B(KEYINPUT90), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n401_), .B(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n395_), .A2(new_n397_), .A3(new_n389_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n404_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n405_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(new_n398_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n379_), .A2(new_n382_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(new_n373_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n410_), .A2(new_n251_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n387_), .A2(new_n410_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT12), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT7), .ZN(new_n416_));
  INV_X1    g215(.A(G99gat), .ZN(new_n417_));
  INV_X1    g216(.A(G106gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT66), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G99gat), .A2(G106gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n419_), .A2(KEYINPUT66), .A3(new_n420_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n423_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(G92gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n206_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT8), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G85gat), .A2(G92gat), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT64), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT9), .B1(new_n433_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n435_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT9), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT64), .B(new_n440_), .C1(new_n206_), .C2(new_n432_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n443_), .A2(new_n444_), .A3(G106gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(new_n428_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n431_), .A2(new_n436_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n419_), .A2(new_n426_), .A3(new_n427_), .A4(new_n420_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT65), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n433_), .A2(new_n435_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n434_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n415_), .B1(new_n447_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G64gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(G57gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n204_), .A2(G64gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT11), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT68), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G57gat), .B(G64gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT68), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(KEYINPUT11), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT67), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT11), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n204_), .A2(G64gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n455_), .A2(G57gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n465_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G71gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(G78gat), .ZN(new_n470_));
  INV_X1    g269(.A(G78gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G71gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n464_), .B1(new_n468_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT11), .B1(new_n456_), .B2(new_n457_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G71gat), .B(G78gat), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n475_), .A2(KEYINPUT67), .A3(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n463_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT67), .B1(new_n475_), .B2(new_n476_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n473_), .B(new_n464_), .C1(new_n460_), .C2(KEYINPUT11), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n479_), .A2(new_n459_), .A3(new_n462_), .A4(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n478_), .A2(KEYINPUT69), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT69), .B1(new_n478_), .B2(new_n481_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n454_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT70), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT70), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n454_), .B(new_n486_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n447_), .A2(new_n453_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n478_), .A2(new_n481_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n415_), .ZN(new_n491_));
  AND2_X1   g290(.A1(G230gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n488_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n489_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n485_), .A2(new_n487_), .A3(new_n491_), .A4(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n494_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n490_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n492_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n484_), .A2(KEYINPUT70), .B1(new_n415_), .B2(new_n490_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n502_), .A2(KEYINPUT71), .A3(new_n487_), .A4(new_n495_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n498_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G120gat), .B(G148gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(new_n293_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT5), .B(G176gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n498_), .A2(new_n501_), .A3(new_n503_), .A4(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(KEYINPUT13), .A3(new_n511_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G8gat), .ZN(new_n517_));
  INV_X1    g316(.A(G1gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT79), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT79), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(G1gat), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n517_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT14), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n518_), .B(new_n519_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT79), .B(G1gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(new_n527_), .B2(new_n517_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n518_), .B1(new_n528_), .B2(new_n519_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n517_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n520_), .A2(new_n522_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n524_), .B1(new_n531_), .B2(G8gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n519_), .ZN(new_n533_));
  OAI21_X1  g332(.A(G1gat), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(G8gat), .A3(new_n525_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(G36gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(G29gat), .ZN(new_n538_));
  INV_X1    g337(.A(G29gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G36gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(G50gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G43gat), .ZN(new_n543_));
  INV_X1    g342(.A(G43gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(G50gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n538_), .A2(new_n540_), .A3(new_n543_), .A4(new_n545_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT81), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(KEYINPUT81), .A3(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT82), .B1(new_n536_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT82), .ZN(new_n556_));
  AOI211_X1 g355(.A(new_n556_), .B(new_n553_), .C1(new_n530_), .C2(new_n535_), .ZN(new_n557_));
  OAI22_X1  g356(.A1(new_n555_), .A2(new_n557_), .B1(new_n536_), .B2(new_n554_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n541_), .A2(new_n546_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n538_), .A2(new_n540_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT73), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT73), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n547_), .A2(new_n565_), .A3(new_n548_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n564_), .A2(new_n566_), .A3(KEYINPUT15), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT15), .B1(new_n564_), .B2(new_n566_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT83), .B1(new_n569_), .B2(new_n536_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT15), .ZN(new_n571_));
  INV_X1    g370(.A(new_n566_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n565_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n564_), .A2(new_n566_), .A3(KEYINPUT15), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT83), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n535_), .A4(new_n530_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n570_), .A2(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n534_), .A2(G8gat), .A3(new_n525_), .ZN(new_n580_));
  AOI21_X1  g379(.A(G8gat), .B1(new_n534_), .B2(new_n525_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n554_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n556_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n536_), .A2(KEYINPUT82), .A3(new_n554_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n579_), .A2(new_n585_), .A3(new_n559_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT84), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G169gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(new_n295_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT85), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n561_), .A2(new_n586_), .B1(new_n587_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n561_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n591_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n590_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n593_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n516_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n414_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G134gat), .ZN(new_n605_));
  INV_X1    g404(.A(G162gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT75), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT72), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n493_), .A2(new_n549_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n493_), .A2(new_n569_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n616_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n619_), .A2(new_n616_), .A3(new_n620_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n607_), .B(new_n608_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT76), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n623_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n625_), .A2(new_n626_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT37), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n622_), .A2(new_n621_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n624_), .B1(new_n630_), .B2(KEYINPUT77), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n622_), .A2(new_n632_), .A3(new_n621_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n623_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n629_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G127gat), .B(G155gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT16), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(G183gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(G211gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT17), .Z(new_n643_));
  NAND2_X1  g442(.A1(G231gat), .A2(G233gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT80), .Z(new_n645_));
  NAND3_X1  g444(.A1(new_n530_), .A2(new_n535_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n489_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n648_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n494_), .A3(new_n646_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n643_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n650_), .B(new_n646_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n482_), .A2(new_n483_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n654_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n653_), .A2(new_n655_), .A3(KEYINPUT17), .A4(new_n642_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n638_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n601_), .A2(new_n658_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n659_), .A2(KEYINPUT105), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(KEYINPUT105), .ZN(new_n661_));
  INV_X1    g460(.A(new_n251_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n531_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT106), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n660_), .A2(new_n666_), .A3(new_n661_), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT38), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n634_), .A2(new_n623_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n414_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n600_), .A2(new_n657_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n675_), .B2(new_n662_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n665_), .A2(KEYINPUT38), .A3(new_n667_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n670_), .A2(new_n676_), .A3(new_n677_), .ZN(G1324gat));
  NAND4_X1  g477(.A1(new_n660_), .A2(new_n517_), .A3(new_n411_), .A4(new_n661_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n387_), .A2(new_n410_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n413_), .A2(new_n412_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n682_), .A2(new_n671_), .A3(new_n411_), .A4(new_n674_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT107), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT39), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n517_), .B1(new_n683_), .B2(KEYINPUT107), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n679_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1325gat));
  AND2_X1   g490(.A1(new_n660_), .A2(new_n661_), .ZN(new_n692_));
  INV_X1    g491(.A(G15gat), .ZN(new_n693_));
  INV_X1    g492(.A(new_n410_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G15gat), .B1(new_n675_), .B2(new_n410_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n698_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n695_), .A2(new_n699_), .A3(new_n700_), .ZN(G1326gat));
  INV_X1    g500(.A(G22gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n692_), .A2(new_n702_), .A3(new_n373_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G22gat), .B1(new_n675_), .B2(new_n374_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT42), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1327gat));
  INV_X1    g505(.A(new_n657_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n671_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n601_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G29gat), .B1(new_n710_), .B2(new_n251_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n599_), .A2(new_n657_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n414_), .B2(new_n637_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  AOI22_X1  g513(.A1(new_n374_), .A2(new_n346_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n694_), .B1(new_n715_), .B2(new_n386_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n413_), .A2(new_n412_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n714_), .B(new_n638_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n712_), .B1(new_n713_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT44), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n721_), .A2(new_n539_), .A3(new_n662_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n719_), .A2(KEYINPUT44), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n711_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(new_n411_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(G36gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n710_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT45), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n720_), .A2(new_n411_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n719_), .A2(KEYINPUT44), .ZN(new_n730_));
  OAI21_X1  g529(.A(G36gat), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n728_), .A2(new_n731_), .A3(KEYINPUT46), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1329gat));
  OAI21_X1  g535(.A(new_n544_), .B1(new_n709_), .B2(new_n410_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n720_), .A2(G43gat), .A3(new_n694_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(new_n730_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g539(.A(G50gat), .B1(new_n710_), .B2(new_n373_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n721_), .A2(new_n542_), .A3(new_n374_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n723_), .ZN(G1331gat));
  AND2_X1   g542(.A1(new_n514_), .A2(new_n515_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n414_), .A2(new_n597_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n658_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n204_), .B1(new_n746_), .B2(new_n662_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n597_), .A2(new_n657_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n673_), .A2(new_n516_), .A3(new_n748_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n749_), .A2(new_n204_), .A3(new_n662_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n750_), .B2(KEYINPUT109), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(KEYINPUT109), .B2(new_n750_), .ZN(G1332gat));
  OAI21_X1  g551(.A(G64gat), .B1(new_n749_), .B2(new_n725_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT48), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n411_), .A2(new_n455_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n746_), .B2(new_n755_), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n749_), .B2(new_n410_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT49), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n694_), .A2(new_n469_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n746_), .B2(new_n759_), .ZN(G1334gat));
  OAI21_X1  g559(.A(G78gat), .B1(new_n749_), .B2(new_n374_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT50), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n373_), .A2(new_n471_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n746_), .B2(new_n763_), .ZN(G1335gat));
  NAND2_X1  g563(.A1(new_n745_), .A2(new_n708_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n206_), .B1(new_n765_), .B2(new_n662_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT110), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n516_), .A2(new_n657_), .A3(new_n598_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n713_), .B2(new_n718_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n770_), .A2(new_n206_), .A3(new_n662_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n767_), .A2(new_n771_), .ZN(G1336gat));
  OAI21_X1  g571(.A(G92gat), .B1(new_n770_), .B2(new_n725_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n765_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n432_), .A3(new_n411_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1337gat));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT112), .B1(new_n777_), .B2(KEYINPUT111), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(KEYINPUT112), .B2(new_n777_), .ZN(new_n779_));
  NOR4_X1   g578(.A1(new_n765_), .A2(new_n444_), .A3(new_n443_), .A4(new_n410_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n417_), .B1(new_n769_), .B2(new_n694_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  MUX2_X1   g581(.A(new_n778_), .B(new_n779_), .S(new_n782_), .Z(G1338gat));
  AOI21_X1  g582(.A(new_n418_), .B1(new_n769_), .B2(new_n373_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n784_), .B2(KEYINPUT113), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n374_), .B(new_n768_), .C1(new_n713_), .C2(new_n718_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n418_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n774_), .A2(new_n418_), .A3(new_n373_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n786_), .B2(new_n418_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(KEYINPUT52), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT53), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n784_), .A2(KEYINPUT113), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n791_), .A3(KEYINPUT52), .ZN(new_n795_));
  OR3_X1    g594(.A1(new_n784_), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .A4(new_n790_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n793_), .A2(new_n798_), .ZN(G1339gat));
  NAND2_X1  g598(.A1(new_n725_), .A2(new_n251_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n410_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n496_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n485_), .A2(new_n499_), .A3(new_n487_), .A4(new_n491_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n802_), .A2(KEYINPUT55), .B1(new_n492_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n498_), .A2(new_n805_), .A3(new_n503_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT56), .A3(new_n509_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT118), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n498_), .A2(new_n805_), .A3(new_n503_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n803_), .A2(new_n492_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n805_), .B2(new_n496_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n810_), .B(new_n509_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT117), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n807_), .A2(new_n810_), .A3(new_n509_), .A4(new_n816_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n809_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n593_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n560_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n558_), .A2(new_n560_), .B1(new_n822_), .B2(new_n579_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT85), .B1(new_n823_), .B2(new_n587_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n821_), .B(new_n511_), .C1(new_n824_), .C2(new_n590_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(KEYINPUT116), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n597_), .B2(new_n511_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n820_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n558_), .A2(new_n559_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n596_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(KEYINPUT119), .A3(new_n596_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n579_), .A2(new_n585_), .A3(new_n560_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n823_), .A2(new_n590_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n512_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n830_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n671_), .A2(KEYINPUT57), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n837_), .A2(new_n838_), .A3(new_n511_), .ZN(new_n844_));
  AOI211_X1 g643(.A(new_n815_), .B(new_n508_), .C1(new_n804_), .C2(new_n806_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT56), .B1(new_n807_), .B2(new_n509_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n844_), .B(KEYINPUT58), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n846_), .B2(new_n845_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n637_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n841_), .A2(new_n843_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n820_), .A2(new_n829_), .B1(new_n512_), .B2(new_n839_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n672_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n707_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n514_), .A2(new_n748_), .A3(new_n515_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT114), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n856_), .A2(KEYINPUT114), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n637_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n744_), .A2(new_n864_), .A3(new_n748_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n857_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n637_), .A3(new_n861_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n863_), .A2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n374_), .B(new_n801_), .C1(new_n855_), .C2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT59), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n841_), .B2(new_n671_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n848_), .A2(new_n849_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n638_), .A3(new_n847_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n853_), .B2(new_n842_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n657_), .B1(new_n871_), .B2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n861_), .B1(new_n866_), .B2(new_n637_), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n638_), .B(new_n862_), .C1(new_n865_), .C2(new_n857_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(new_n374_), .A4(new_n801_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n870_), .A2(new_n597_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G113gat), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n598_), .A2(G113gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n869_), .B2(new_n884_), .ZN(G1340gat));
  NAND3_X1  g684(.A1(new_n870_), .A2(new_n516_), .A3(new_n881_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n870_), .A2(KEYINPUT120), .A3(new_n516_), .A4(new_n881_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(G120gat), .A3(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n855_), .A2(new_n868_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n373_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n744_), .A2(G120gat), .ZN(new_n893_));
  MUX2_X1   g692(.A(new_n893_), .B(G120gat), .S(KEYINPUT60), .Z(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n801_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n890_), .A2(new_n895_), .ZN(G1341gat));
  NAND3_X1  g695(.A1(new_n870_), .A2(new_n707_), .A3(new_n881_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G127gat), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n657_), .A2(G127gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n869_), .B2(new_n899_), .ZN(G1342gat));
  NAND3_X1  g699(.A1(new_n870_), .A2(new_n638_), .A3(new_n881_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G134gat), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n671_), .A2(G134gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n869_), .B2(new_n903_), .ZN(G1343gat));
  NAND2_X1  g703(.A1(new_n410_), .A2(new_n373_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n800_), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT121), .Z(new_n907_));
  NAND2_X1  g706(.A1(new_n879_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n598_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT122), .B(G141gat), .Z(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1344gat));
  NOR2_X1   g710(.A1(new_n908_), .A2(new_n744_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n213_), .ZN(G1345gat));
  NOR2_X1   g712(.A1(new_n908_), .A2(new_n657_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT61), .B(G155gat), .Z(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1346gat));
  NOR3_X1   g715(.A1(new_n908_), .A2(new_n606_), .A3(new_n637_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n606_), .B1(new_n908_), .B2(new_n671_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n919_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n917_), .B1(new_n920_), .B2(new_n921_), .ZN(G1347gat));
  NAND2_X1  g721(.A1(new_n413_), .A2(new_n411_), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT124), .Z(new_n924_));
  NAND3_X1  g723(.A1(new_n879_), .A2(new_n374_), .A3(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925_), .B2(new_n598_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n892_), .A2(new_n280_), .A3(new_n597_), .A4(new_n924_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n927_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n928_), .A2(new_n929_), .A3(new_n930_), .ZN(G1348gat));
  NOR2_X1   g730(.A1(new_n925_), .A2(new_n744_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n281_), .ZN(G1349gat));
  INV_X1    g732(.A(new_n265_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n892_), .A2(new_n707_), .A3(new_n934_), .A4(new_n924_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n269_), .B1(new_n925_), .B2(new_n657_), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n925_), .B2(new_n637_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n672_), .A2(new_n266_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n925_), .B2(new_n942_), .ZN(G1351gat));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n905_), .A2(new_n725_), .A3(new_n251_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n879_), .B2(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n945_), .ZN(new_n947_));
  AOI211_X1 g746(.A(KEYINPUT126), .B(new_n947_), .C1(new_n875_), .C2(new_n878_), .ZN(new_n948_));
  OAI211_X1 g747(.A(G197gat), .B(new_n597_), .C1(new_n946_), .C2(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  OAI21_X1  g750(.A(KEYINPUT126), .B1(new_n891_), .B2(new_n947_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n879_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n954_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n597_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n597_), .B1(new_n946_), .B2(new_n948_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n295_), .ZN(new_n957_));
  AND3_X1   g756(.A1(new_n951_), .A2(new_n955_), .A3(new_n957_), .ZN(G1352gat));
  NOR2_X1   g757(.A1(new_n946_), .A2(new_n948_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n959_), .A2(new_n293_), .A3(new_n744_), .ZN(new_n960_));
  AOI21_X1  g759(.A(G204gat), .B1(new_n954_), .B2(new_n516_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1353gat));
  OR2_X1    g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n963_), .B1(new_n954_), .B2(new_n707_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n959_), .A2(new_n657_), .ZN(new_n965_));
  XOR2_X1   g764(.A(KEYINPUT63), .B(G211gat), .Z(new_n966_));
  AOI21_X1  g765(.A(new_n964_), .B1(new_n965_), .B2(new_n966_), .ZN(G1354gat));
  OR3_X1    g766(.A1(new_n959_), .A2(G218gat), .A3(new_n671_), .ZN(new_n968_));
  OAI21_X1  g767(.A(G218gat), .B1(new_n959_), .B2(new_n637_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1355gat));
endmodule


