//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n204_));
  AND2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n211_), .B(new_n212_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT83), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n214_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n213_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n208_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n207_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n209_), .B1(new_n205_), .B2(KEYINPUT1), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n204_), .B1(new_n220_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n214_), .B(KEYINPUT83), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(KEYINPUT2), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n207_), .B1(new_n228_), .B2(new_n215_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT84), .A3(new_n224_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n226_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT28), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G228gat), .A2(G233gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT86), .Z(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n226_), .A2(new_n230_), .A3(KEYINPUT29), .ZN(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(G204gat), .ZN(new_n240_));
  INV_X1    g039(.A(G204gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(G197gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT21), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT87), .B1(new_n239_), .B2(G204gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT87), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(new_n241_), .A3(G197gat), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n245_), .B(new_n247_), .C1(G197gat), .C2(new_n241_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n243_), .B(new_n244_), .C1(new_n248_), .C2(KEYINPUT21), .ZN(new_n249_));
  INV_X1    g048(.A(new_n244_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(KEYINPUT21), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n237_), .B1(new_n238_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G78gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n220_), .A2(new_n225_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n237_), .B(new_n252_), .C1(new_n255_), .C2(new_n232_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n253_), .A2(new_n254_), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n254_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G106gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT85), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(G106gat), .A3(new_n259_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n234_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT85), .ZN(new_n265_));
  INV_X1    g064(.A(new_n259_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n253_), .A2(new_n257_), .A3(new_n254_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n261_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AND4_X1   g067(.A1(new_n265_), .A2(new_n268_), .A3(new_n263_), .A4(new_n234_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n203_), .B1(new_n264_), .B2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n234_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n262_), .A2(new_n234_), .A3(new_n263_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n202_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(G169gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(G183gat), .A3(G190gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G183gat), .ZN(new_n283_));
  INV_X1    g082(.A(G190gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT23), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n278_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT79), .ZN(new_n290_));
  INV_X1    g089(.A(G169gat), .ZN(new_n291_));
  INV_X1    g090(.A(G176gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT24), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G190gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT25), .B(G183gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT24), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n285_), .A2(new_n280_), .B1(new_n298_), .B2(new_n289_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n294_), .B(new_n297_), .C1(KEYINPUT90), .C2(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(KEYINPUT90), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n288_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT20), .B1(new_n302_), .B2(new_n252_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n252_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT78), .B(G183gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n284_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n285_), .A2(new_n280_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n278_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n282_), .A2(new_n285_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n295_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n290_), .A2(new_n298_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n294_), .A2(new_n313_), .A3(new_n317_), .A4(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n307_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n303_), .A2(new_n306_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n302_), .A2(new_n252_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n307_), .A2(new_n319_), .A3(new_n312_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT89), .B1(new_n323_), .B2(KEYINPUT20), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n306_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G64gat), .B(G92gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT92), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  AND3_X1   g132(.A1(new_n321_), .A2(new_n327_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n321_), .A2(new_n327_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n333_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT93), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n321_), .A2(new_n327_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(KEYINPUT93), .A3(new_n333_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n325_), .A2(new_n326_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n303_), .A2(new_n320_), .ZN(new_n345_));
  MUX2_X1   g144(.A(new_n344_), .B(new_n345_), .S(new_n306_), .Z(new_n346_));
  OAI211_X1 g145(.A(KEYINPUT27), .B(new_n335_), .C1(new_n346_), .C2(new_n333_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n319_), .A2(new_n312_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT30), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT81), .B(G43gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G15gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(G71gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G113gat), .B(G120gat), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n359_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(KEYINPUT82), .A3(new_n361_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT31), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G99gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n352_), .A2(new_n355_), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n357_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n357_), .B2(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n226_), .A2(new_n366_), .A3(new_n230_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n255_), .A2(new_n362_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n374_), .A2(new_n375_), .A3(KEYINPUT4), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n226_), .A2(new_n366_), .A3(new_n230_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT94), .B1(new_n376_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G85gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT0), .B(G57gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n384_), .B(new_n385_), .Z(new_n386_));
  NAND3_X1  g185(.A1(new_n374_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n374_), .A2(new_n375_), .A3(KEYINPUT4), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT94), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(new_n380_), .A4(new_n378_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n382_), .A2(new_n386_), .A3(new_n387_), .A4(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n391_), .A2(KEYINPUT96), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(KEYINPUT96), .ZN(new_n393_));
  INV_X1    g192(.A(new_n386_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n382_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n387_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n392_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n398_));
  NOR4_X1   g197(.A1(new_n276_), .A2(new_n348_), .A3(new_n373_), .A4(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT97), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n339_), .A2(new_n341_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n390_), .A2(new_n387_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n402_), .A2(KEYINPUT33), .A3(new_n386_), .A4(new_n382_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n374_), .A2(new_n375_), .A3(new_n380_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n404_), .A2(new_n394_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(KEYINPUT95), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(KEYINPUT95), .A3(new_n394_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n388_), .A2(new_n379_), .A3(new_n378_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n391_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n403_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT32), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n336_), .B1(new_n414_), .B2(new_n337_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n337_), .A2(new_n414_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n306_), .B1(new_n303_), .B2(new_n320_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n416_), .B(new_n417_), .C1(new_n344_), .C2(new_n306_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n401_), .A2(new_n413_), .B1(new_n398_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n400_), .B1(new_n276_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n397_), .B1(KEYINPUT96), .B2(new_n391_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n393_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n333_), .B1(new_n321_), .B2(new_n327_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n334_), .A2(new_n425_), .A3(KEYINPUT93), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n340_), .A2(KEYINPUT93), .A3(new_n333_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n428_), .B2(new_n412_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n429_), .A2(KEYINPUT97), .A3(new_n275_), .A4(new_n270_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n422_), .A2(new_n423_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n343_), .A2(new_n347_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n276_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n421_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n399_), .B1(new_n434_), .B2(new_n373_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT74), .B(G1gat), .ZN(new_n436_));
  INV_X1    g235(.A(G8gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT14), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G1gat), .B(G8gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G29gat), .B(G36gat), .Z(new_n443_));
  XOR2_X1   g242(.A(G43gat), .B(G50gat), .Z(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  XNOR2_X1  g244(.A(new_n442_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G229gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT76), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT76), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n446_), .A2(new_n451_), .A3(new_n448_), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n445_), .B(KEYINPUT15), .Z(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n442_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n442_), .A2(new_n445_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n455_), .A2(new_n447_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n450_), .A2(new_n452_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G113gat), .B(G141gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT77), .ZN(new_n459_));
  XOR2_X1   g258(.A(G169gat), .B(G197gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(new_n462_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n435_), .A2(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n468_), .A2(KEYINPUT64), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT64), .B1(new_n468_), .B2(new_n469_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n261_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT6), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G85gat), .A2(G92gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(new_n476_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT9), .B1(new_n479_), .B2(KEYINPUT65), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT9), .ZN(new_n482_));
  NOR4_X1   g281(.A1(new_n478_), .A2(new_n476_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n477_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT66), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT66), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n486_), .B(new_n477_), .C1(new_n480_), .C2(new_n483_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n475_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT69), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n479_), .A2(KEYINPUT8), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n473_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT67), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT7), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n495_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n492_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT68), .B(new_n496_), .C1(new_n497_), .C2(new_n495_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n490_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n474_), .B(new_n496_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT8), .B1(new_n503_), .B2(new_n479_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n489_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT67), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n495_), .B1(new_n494_), .B2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n494_), .A2(new_n495_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n499_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(new_n474_), .A3(new_n501_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n490_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n479_), .B1(new_n498_), .B2(new_n492_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n513_), .A2(KEYINPUT69), .A3(new_n516_), .ZN(new_n517_));
  AOI211_X1 g316(.A(KEYINPUT70), .B(new_n488_), .C1(new_n505_), .C2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT70), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n505_), .A2(new_n517_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n488_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n453_), .B1(new_n518_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT34), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n488_), .A2(new_n504_), .A3(new_n502_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n445_), .ZN(new_n531_));
  AOI211_X1 g330(.A(new_n528_), .B(new_n529_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n527_), .A3(new_n526_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n527_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n523_), .A2(new_n535_), .A3(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G190gat), .B(G218gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G134gat), .B(G162gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(KEYINPUT36), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n540_), .B(KEYINPUT36), .Z(new_n545_));
  NAND3_X1  g344(.A1(new_n534_), .A2(new_n536_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT37), .B1(new_n542_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G57gat), .B(G64gat), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT11), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(KEYINPUT11), .ZN(new_n553_));
  XOR2_X1   g352(.A(G71gat), .B(G78gat), .Z(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n553_), .A2(new_n554_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n442_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G127gat), .B(G155gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT17), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(KEYINPUT17), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n560_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n566_), .B2(new_n560_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n550_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n557_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT12), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n518_), .B2(new_n522_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n530_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n572_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n530_), .B2(new_n557_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n575_), .A2(new_n579_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n530_), .A2(new_n557_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n581_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G120gat), .B(G148gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n583_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT71), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AOI211_X1 g394(.A(KEYINPUT71), .B(new_n591_), .C1(new_n583_), .C2(new_n586_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n597_));
  OAI22_X1  g396(.A1(new_n595_), .A2(new_n596_), .B1(KEYINPUT72), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n583_), .A2(new_n586_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n590_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(KEYINPUT71), .A3(new_n592_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n596_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n571_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n467_), .A2(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n609_), .A2(KEYINPUT99), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(KEYINPUT99), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n610_), .A2(new_n398_), .A3(new_n436_), .A4(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n542_), .A2(new_n548_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n435_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n606_), .A2(new_n465_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(new_n569_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(new_n431_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n612_), .A2(new_n613_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n614_), .A2(new_n620_), .A3(new_n621_), .ZN(G1324gat));
  NAND3_X1  g421(.A1(new_n616_), .A2(new_n348_), .A3(new_n618_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(G8gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT39), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n610_), .A2(new_n437_), .A3(new_n348_), .A4(new_n611_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(G1325gat));
  OAI21_X1  g428(.A(G15gat), .B1(new_n619_), .B2(new_n373_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n609_), .A2(G15gat), .A3(new_n373_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(new_n276_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G22gat), .B1(new_n619_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT42), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n634_), .A2(G22gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n609_), .B2(new_n637_), .ZN(G1327gat));
  INV_X1    g437(.A(new_n615_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n607_), .A2(new_n570_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n467_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n398_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT101), .B1(new_n435_), .B2(new_n550_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT101), .B(KEYINPUT43), .C1(new_n435_), .C2(new_n550_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n617_), .A2(new_n570_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT44), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651_));
  INV_X1    g450(.A(new_n649_), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n651_), .B(new_n652_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n398_), .A2(G29gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n643_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(G36gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n348_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n641_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n348_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n650_), .A2(new_n653_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n663_), .B2(new_n657_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n661_), .B(new_n665_), .C1(new_n663_), .C2(new_n657_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  INV_X1    g468(.A(new_n550_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n373_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n412_), .B1(new_n341_), .B2(new_n339_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n391_), .A2(KEYINPUT96), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n386_), .B1(new_n402_), .B2(new_n382_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI22_X1  g474(.A1(new_n675_), .A2(new_n393_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n270_), .B(new_n275_), .C1(new_n672_), .C2(new_n676_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n677_), .A2(new_n400_), .B1(new_n276_), .B2(new_n432_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n671_), .B1(new_n678_), .B2(new_n430_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n670_), .B1(new_n679_), .B2(new_n399_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT43), .B1(new_n680_), .B2(KEYINPUT101), .ZN(new_n681_));
  INV_X1    g480(.A(new_n647_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n651_), .B1(new_n683_), .B2(new_n652_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n649_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n684_), .A2(G43gat), .A3(new_n671_), .A4(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G43gat), .B1(new_n642_), .B2(new_n671_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n684_), .A2(new_n276_), .A3(new_n685_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G50gat), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n641_), .A2(G50gat), .A3(new_n634_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n691_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT104), .B(new_n694_), .C1(new_n692_), .C2(G50gat), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1331gat));
  NOR2_X1   g497(.A1(new_n435_), .A2(new_n465_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n571_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n607_), .A3(new_n700_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT105), .Z(new_n702_));
  INV_X1    g501(.A(G57gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n398_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n606_), .A2(new_n465_), .A3(new_n569_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n616_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n431_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n702_), .A2(new_n709_), .A3(new_n348_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G64gat), .B1(new_n706_), .B2(new_n662_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1333gat));
  NOR2_X1   g512(.A1(new_n373_), .A2(G71gat), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT106), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n702_), .A2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G71gat), .B1(new_n706_), .B2(new_n373_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT49), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1334gat));
  NAND2_X1  g518(.A1(new_n276_), .A2(new_n254_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT107), .Z(new_n721_));
  NAND2_X1  g520(.A1(new_n702_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n616_), .A2(new_n276_), .A3(new_n705_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G78gat), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n465_), .A2(new_n570_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n607_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n648_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n431_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n699_), .A2(new_n607_), .A3(new_n569_), .A4(new_n615_), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n734_), .A2(G85gat), .A3(new_n431_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1336gat));
  OAI21_X1  g535(.A(G92gat), .B1(new_n732_), .B2(new_n662_), .ZN(new_n737_));
  OR3_X1    g536(.A1(new_n734_), .A2(G92gat), .A3(new_n662_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1337gat));
  NAND3_X1  g538(.A1(new_n648_), .A2(new_n671_), .A3(new_n731_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(G99gat), .ZN(new_n741_));
  INV_X1    g540(.A(new_n734_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n470_), .A2(new_n471_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(new_n671_), .A3(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n741_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(G1338gat));
  OAI211_X1 g546(.A(new_n276_), .B(new_n731_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n748_), .A2(KEYINPUT109), .A3(G106gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT109), .B1(new_n748_), .B2(G106gat), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n634_), .B(new_n730_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n753_), .B(new_n751_), .C1(new_n754_), .C2(new_n261_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n742_), .A2(new_n261_), .A3(new_n276_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT53), .B1(new_n752_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n753_), .B1(new_n754_), .B2(new_n261_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n748_), .A2(KEYINPUT109), .A3(G106gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(KEYINPUT52), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n755_), .A4(new_n756_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(G113gat), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n454_), .A2(new_n455_), .A3(new_n448_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n462_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n457_), .A2(new_n462_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n592_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n575_), .A2(new_n584_), .A3(new_n579_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n581_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n583_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n575_), .A2(new_n579_), .A3(KEYINPUT55), .A4(new_n582_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n590_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n590_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n771_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n767_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n771_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n590_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n590_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(KEYINPUT114), .A3(KEYINPUT58), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n784_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n766_), .B1(new_n790_), .B2(new_n670_), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT115), .B(new_n550_), .C1(new_n784_), .C2(new_n789_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n465_), .A2(new_n592_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n601_), .A2(new_n602_), .A3(new_n770_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n615_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT57), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT112), .B(KEYINPUT57), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n797_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n801_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n601_), .A2(new_n602_), .A3(new_n770_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n780_), .A2(new_n781_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n794_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT113), .B(new_n803_), .C1(new_n806_), .C2(new_n615_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n799_), .B1(new_n802_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n570_), .B1(new_n793_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n465_), .A2(new_n569_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n601_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n597_), .A2(KEYINPUT72), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n810_), .B(new_n811_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n550_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n810_), .B1(new_n606_), .B2(new_n811_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT54), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n811_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT110), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n550_), .A4(new_n815_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT116), .B1(new_n809_), .B2(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n788_), .A2(KEYINPUT114), .A3(KEYINPUT58), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT58), .B1(new_n788_), .B2(KEYINPUT114), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n670_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT115), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n802_), .A2(new_n807_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n790_), .A2(new_n766_), .A3(new_n670_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n828_), .A2(new_n829_), .A3(new_n798_), .A4(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n569_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833_));
  INV_X1    g632(.A(new_n823_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  NOR4_X1   g634(.A1(new_n276_), .A2(new_n348_), .A3(new_n373_), .A4(new_n431_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n824_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n765_), .B1(new_n837_), .B2(new_n466_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT117), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n840_), .B(new_n765_), .C1(new_n837_), .C2(new_n466_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n827_), .B(new_n798_), .C1(new_n797_), .C2(new_n801_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n569_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n834_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n836_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n837_), .B2(KEYINPUT59), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n466_), .A2(new_n765_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n839_), .A2(new_n841_), .B1(new_n847_), .B2(new_n848_), .ZN(G1340gat));
  AOI211_X1 g648(.A(new_n606_), .B(new_n846_), .C1(new_n837_), .C2(KEYINPUT59), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n606_), .B2(KEYINPUT60), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n851_), .A2(KEYINPUT60), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n850_), .A2(new_n851_), .B1(new_n837_), .B2(new_n854_), .ZN(G1341gat));
  AOI211_X1 g654(.A(new_n569_), .B(new_n846_), .C1(new_n837_), .C2(KEYINPUT59), .ZN(new_n856_));
  INV_X1    g655(.A(G127gat), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n570_), .A2(new_n857_), .ZN(new_n858_));
  OAI22_X1  g657(.A1(new_n856_), .A2(new_n857_), .B1(new_n837_), .B2(new_n858_), .ZN(G1342gat));
  AOI211_X1 g658(.A(new_n550_), .B(new_n846_), .C1(new_n837_), .C2(KEYINPUT59), .ZN(new_n860_));
  INV_X1    g659(.A(G134gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n615_), .A2(new_n861_), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n860_), .A2(new_n861_), .B1(new_n837_), .B2(new_n862_), .ZN(G1343gat));
  XNOR2_X1  g662(.A(KEYINPUT119), .B(G141gat), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n276_), .A2(new_n662_), .A3(new_n398_), .A4(new_n373_), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT118), .Z(new_n867_));
  NAND4_X1  g666(.A1(new_n824_), .A2(new_n465_), .A3(new_n835_), .A4(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n865_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n864_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(G1344gat));
  AOI21_X1  g674(.A(new_n833_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n876_));
  AOI211_X1 g675(.A(KEYINPUT116), .B(new_n823_), .C1(new_n831_), .C2(new_n569_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n607_), .A3(new_n867_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n878_), .A2(new_n881_), .A3(new_n570_), .A4(new_n867_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n824_), .A2(new_n570_), .A3(new_n835_), .A4(new_n867_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT121), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n882_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1346gat));
  NAND3_X1  g687(.A1(new_n878_), .A2(new_n670_), .A3(new_n867_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G162gat), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n639_), .A2(G162gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n878_), .A2(new_n867_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1347gat));
  NAND3_X1  g692(.A1(new_n671_), .A2(new_n348_), .A3(new_n431_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT122), .Z(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n276_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n844_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n465_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  AND4_X1   g700(.A1(KEYINPUT123), .A2(new_n900_), .A3(new_n901_), .A4(G169gat), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n291_), .B1(new_n903_), .B2(KEYINPUT62), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n900_), .A2(new_n904_), .B1(KEYINPUT123), .B2(new_n901_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT22), .B(G169gat), .Z(new_n906_));
  OAI22_X1  g705(.A1(new_n902_), .A2(new_n905_), .B1(new_n900_), .B2(new_n906_), .ZN(G1348gat));
  NOR3_X1   g706(.A1(new_n896_), .A2(new_n292_), .A3(new_n606_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n878_), .A2(new_n634_), .A3(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n292_), .B1(new_n898_), .B2(new_n606_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n909_), .A2(KEYINPUT124), .A3(new_n910_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1349gat));
  NOR3_X1   g714(.A1(new_n898_), .A2(new_n296_), .A3(new_n569_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n878_), .A2(new_n634_), .A3(new_n570_), .A4(new_n895_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n308_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n898_), .B2(new_n550_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n615_), .A2(new_n295_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n898_), .B2(new_n920_), .ZN(G1351gat));
  NOR4_X1   g720(.A1(new_n634_), .A2(new_n662_), .A3(new_n398_), .A4(new_n671_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n878_), .A2(new_n465_), .A3(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT125), .B(G197gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n923_), .B2(new_n926_), .ZN(G1352gat));
  NAND3_X1  g726(.A1(new_n878_), .A2(new_n607_), .A3(new_n922_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g728(.A1(new_n824_), .A2(new_n570_), .A3(new_n835_), .A4(new_n922_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT63), .B(G211gat), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n933_));
  INV_X1    g732(.A(G211gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n930_), .A2(KEYINPUT126), .A3(new_n933_), .A4(new_n934_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n932_), .B1(new_n937_), .B2(new_n938_), .ZN(G1354gat));
  NAND3_X1  g738(.A1(new_n878_), .A2(new_n670_), .A3(new_n922_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(G218gat), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n639_), .A2(G218gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n878_), .A2(new_n922_), .A3(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1355gat));
endmodule


