//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT64), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT10), .B(G99gat), .Z(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  OR3_X1    g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT9), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n209_), .A2(new_n212_), .A3(new_n214_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT7), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n209_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n208_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n219_), .B1(new_n224_), .B2(new_n213_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n218_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(KEYINPUT65), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(KEYINPUT65), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G57gat), .B(G64gat), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n232_));
  XOR2_X1   g031(.A(G71gat), .B(G78gat), .Z(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n232_), .A2(new_n233_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT66), .Z(new_n237_));
  NAND3_X1  g036(.A1(new_n228_), .A2(new_n229_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n203_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G120gat), .B(G148gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT5), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G176gat), .B(G204gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n236_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n226_), .A2(KEYINPUT12), .A3(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n238_), .B(new_n248_), .C1(new_n240_), .C2(KEYINPUT12), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n241_), .B(new_n246_), .C1(new_n249_), .C2(new_n203_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT67), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n238_), .A2(new_n248_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n252_), .B(new_n202_), .C1(KEYINPUT12), .C2(new_n240_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n241_), .A4(new_n246_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n241_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n245_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT68), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(KEYINPUT68), .A3(new_n258_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT13), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT13), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n256_), .A2(KEYINPUT68), .A3(new_n258_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n259_), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT73), .B(G1gat), .Z(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT74), .B(G8gat), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT14), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G15gat), .B(G22gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G1gat), .B(G8gat), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G29gat), .B(G36gat), .Z(new_n276_));
  XOR2_X1   g075(.A(G43gat), .B(G50gat), .Z(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT15), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n278_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G229gat), .A2(G233gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n275_), .B(new_n281_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(G229gat), .A3(G233gat), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G113gat), .B(G141gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT78), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT79), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G169gat), .B(G197gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  OR2_X1    g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n288_), .A2(new_n293_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n262_), .A2(new_n265_), .A3(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT87), .B(G43gat), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT81), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT81), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(G169gat), .A3(G176gat), .ZN(new_n303_));
  INV_X1    g102(.A(G169gat), .ZN(new_n304_));
  INV_X1    g103(.A(G176gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n301_), .A2(new_n303_), .A3(new_n306_), .A4(KEYINPUT24), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n306_), .A2(KEYINPUT24), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT80), .ZN(new_n309_));
  INV_X1    g108(.A(G190gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n310_), .B2(KEYINPUT26), .ZN(new_n311_));
  INV_X1    g110(.A(G183gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT25), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G183gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT26), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G190gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n310_), .A2(KEYINPUT26), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n309_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n307_), .B(new_n308_), .C1(new_n316_), .C2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT83), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323_));
  AND2_X1   g122(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n324_));
  NOR2_X1   g123(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n322_), .B(new_n323_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  OR2_X1    g126(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n328_));
  NAND2_X1  g127(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT83), .B1(new_n323_), .B2(KEYINPUT23), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n326_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n301_), .A2(new_n303_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n304_), .A2(KEYINPUT22), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT22), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G169gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n334_), .B1(new_n336_), .B2(G169gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n305_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n333_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n327_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n312_), .A2(new_n310_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n323_), .A2(new_n344_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  OAI22_X1  g145(.A1(new_n321_), .A2(new_n332_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT22), .B(G169gat), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n305_), .B(new_n339_), .C1(new_n350_), .C2(new_n334_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n333_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(KEYINPUT85), .C1(new_n332_), .C2(new_n321_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n349_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n356_), .A2(new_n357_), .A3(G99gat), .ZN(new_n358_));
  INV_X1    g157(.A(G99gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n355_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n306_), .A2(KEYINPUT24), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n311_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n310_), .A2(KEYINPUT26), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n317_), .A2(G190gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT80), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n330_), .A2(new_n331_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n326_), .A4(new_n307_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT85), .B1(new_n368_), .B2(new_n353_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n354_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n360_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n349_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n359_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n299_), .B1(new_n358_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n375_), .B(G15gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G71gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(G99gat), .B1(new_n356_), .B2(new_n357_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n371_), .A2(new_n359_), .A3(new_n372_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(new_n298_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n374_), .A2(new_n377_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n377_), .B1(new_n374_), .B2(new_n380_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT31), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G127gat), .B(G134gat), .Z(new_n386_));
  XOR2_X1   g185(.A(G113gat), .B(G120gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n377_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n378_), .A2(new_n379_), .A3(new_n298_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n298_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT31), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n381_), .A3(new_n382_), .A4(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n385_), .A2(new_n389_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n389_), .B1(new_n385_), .B2(new_n395_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G141gat), .A2(G148gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT89), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(KEYINPUT1), .ZN(new_n403_));
  OR2_X1    g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n403_), .B(new_n404_), .C1(KEYINPUT1), .C2(new_n401_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n402_), .B1(new_n401_), .B2(KEYINPUT1), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n399_), .B(new_n400_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  OR3_X1    g206(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT2), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n400_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n389_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n388_), .A2(new_n407_), .A3(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT98), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n420_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n389_), .A2(new_n415_), .A3(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n422_), .B(new_n424_), .C1(new_n418_), .C2(new_n423_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT98), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n428_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT101), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n421_), .A2(new_n425_), .A3(new_n433_), .A4(new_n427_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n428_), .A2(KEYINPUT101), .A3(new_n434_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT103), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n415_), .A2(KEYINPUT29), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(KEYINPUT90), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT21), .ZN(new_n446_));
  INV_X1    g245(.A(G204gat), .ZN(new_n447_));
  INV_X1    g246(.A(G197gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT92), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G197gat), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n447_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G197gat), .A2(G204gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n446_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G218gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(G211gat), .ZN(new_n456_));
  INV_X1    g255(.A(G211gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G218gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n449_), .A2(new_n451_), .A3(new_n447_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n446_), .B1(G197gat), .B2(G204gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n449_), .A2(new_n451_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n453_), .B1(new_n463_), .B2(G204gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n446_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n454_), .A2(new_n462_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT91), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n443_), .B1(new_n445_), .B2(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(KEYINPUT91), .A2(G228gat), .A3(G233gat), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n444_), .B(new_n467_), .C1(KEYINPUT90), .C2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G78gat), .B(G106gat), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n469_), .A2(new_n475_), .A3(new_n471_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n415_), .A2(KEYINPUT29), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n478_), .A2(KEYINPUT28), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(KEYINPUT28), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G22gat), .B(G50gat), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n481_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n478_), .A2(KEYINPUT28), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(KEYINPUT28), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n477_), .B1(new_n482_), .B2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n482_), .A2(new_n486_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT27), .ZN(new_n491_));
  XOR2_X1   g290(.A(G8gat), .B(G36gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G64gat), .B(G92gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n349_), .A2(new_n354_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n467_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT95), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G226gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT19), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n343_), .B(new_n326_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n336_), .A2(G169gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n304_), .A2(KEYINPUT22), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT94), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n335_), .A2(new_n337_), .A3(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n305_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n503_), .A2(new_n509_), .A3(new_n333_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n363_), .A2(new_n364_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n313_), .A2(new_n315_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n361_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n300_), .A2(KEYINPUT24), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT93), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT93), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n300_), .A2(new_n516_), .A3(KEYINPUT24), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n306_), .A3(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n342_), .A2(new_n345_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n513_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n466_), .A2(new_n510_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT20), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n498_), .A2(new_n499_), .A3(new_n502_), .A4(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n349_), .A2(new_n354_), .A3(new_n466_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT20), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n510_), .A2(new_n520_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n527_), .B2(new_n467_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n501_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n524_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n522_), .B1(new_n497_), .B2(new_n467_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n499_), .B1(new_n532_), .B2(new_n502_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n525_), .A2(new_n502_), .A3(new_n528_), .ZN(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT100), .B(new_n535_), .C1(new_n532_), .C2(new_n502_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n496_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT100), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n466_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n538_), .B(new_n501_), .C1(new_n539_), .C2(new_n522_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n536_), .A2(new_n537_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT102), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n496_), .A2(new_n534_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n536_), .A2(KEYINPUT102), .A3(new_n537_), .A4(new_n540_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n491_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n537_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n498_), .A2(new_n502_), .A3(new_n523_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT95), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n548_), .A2(new_n496_), .A3(new_n524_), .A4(new_n530_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n546_), .A2(new_n491_), .A3(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n442_), .B(new_n490_), .C1(new_n545_), .C2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n541_), .A2(new_n542_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n549_), .A3(new_n544_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(KEYINPUT27), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n490_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT103), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n398_), .A2(new_n441_), .A3(new_n551_), .A4(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(KEYINPUT27), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n546_), .A2(new_n491_), .A3(new_n549_), .ZN(new_n559_));
  AOI211_X1 g358(.A(new_n440_), .B(new_n490_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT99), .ZN(new_n561_));
  INV_X1    g360(.A(new_n437_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT33), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n433_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n424_), .B(new_n420_), .C1(new_n418_), .C2(new_n423_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n561_), .B1(new_n562_), .B2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n563_), .B2(new_n437_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n562_), .A2(new_n561_), .A3(KEYINPUT33), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n568_), .A2(new_n549_), .A3(new_n546_), .A4(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n536_), .A2(KEYINPUT32), .A3(new_n496_), .A4(new_n540_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT32), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n534_), .B1(new_n572_), .B2(new_n537_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n440_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n555_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  OAI22_X1  g374(.A1(new_n560_), .A2(new_n575_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n297_), .B1(new_n557_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n228_), .A2(new_n281_), .A3(new_n229_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n226_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT69), .B1(new_n579_), .B2(new_n279_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n279_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n581_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n578_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT70), .ZN(new_n594_));
  XOR2_X1   g393(.A(G134gat), .B(G162gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n601_));
  INV_X1    g400(.A(new_n592_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(KEYINPUT71), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n596_), .B(KEYINPUT36), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n602_), .B2(KEYINPUT71), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n600_), .B(new_n601_), .C1(new_n603_), .C2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n592_), .A2(new_n604_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT37), .B1(new_n607_), .B2(new_n599_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n275_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n236_), .B(KEYINPUT75), .Z(new_n613_));
  AND2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  XOR2_X1   g414(.A(G127gat), .B(G155gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT16), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n620_));
  NOR4_X1   g419(.A1(new_n614_), .A2(new_n615_), .A3(new_n619_), .A4(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n611_), .B(new_n237_), .Z(new_n622_));
  XOR2_X1   g421(.A(new_n619_), .B(KEYINPUT17), .Z(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n609_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT77), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n577_), .A2(new_n627_), .ZN(new_n628_));
  OR3_X1    g427(.A1(new_n628_), .A2(new_n266_), .A3(new_n441_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT104), .ZN(new_n632_));
  INV_X1    g431(.A(new_n297_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n391_), .A2(new_n392_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT88), .B1(new_n634_), .B2(new_n377_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n394_), .B1(new_n635_), .B2(new_n393_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n395_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n388_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n385_), .A2(new_n389_), .A3(new_n395_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n556_), .A2(new_n638_), .A3(new_n551_), .A4(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n576_), .B1(new_n640_), .B2(new_n440_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n600_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n642_));
  AND4_X1   g441(.A1(new_n633_), .A2(new_n641_), .A3(new_n642_), .A4(new_n625_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n441_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n632_), .B(new_n645_), .C1(new_n630_), .C2(new_n629_), .ZN(G1324gat));
  INV_X1    g445(.A(new_n554_), .ZN(new_n647_));
  OR3_X1    g446(.A1(new_n628_), .A2(new_n267_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(new_n554_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(G8gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n649_), .B2(G8gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g453(.A(new_n398_), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n628_), .A2(G15gat), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G15gat), .B1(new_n644_), .B2(new_n655_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n657_), .A2(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(G1326gat));
  OAI21_X1  g460(.A(G22gat), .B1(new_n644_), .B2(new_n490_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n490_), .A2(G22gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n628_), .B2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n642_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n625_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n633_), .A2(new_n641_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n440_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n297_), .A2(new_n625_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT43), .B(new_n609_), .C1(new_n557_), .C2(new_n576_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  INV_X1    g474(.A(new_n609_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n641_), .B2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n674_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n673_), .B(KEYINPUT44), .C1(new_n674_), .C2(new_n677_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n440_), .A2(G29gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n672_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n647_), .A2(G36gat), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n633_), .A2(new_n641_), .A3(new_n670_), .A4(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n680_), .A2(new_n554_), .A3(new_n681_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(G36gat), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT108), .B(new_n685_), .C1(new_n691_), .C2(KEYINPUT107), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(G36gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n689_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT46), .B1(new_n691_), .B2(KEYINPUT108), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n692_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(G1329gat));
  AND2_X1   g500(.A1(new_n398_), .A2(G43gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n680_), .A2(new_n681_), .A3(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT109), .ZN(new_n704_));
  AOI21_X1  g503(.A(G43gat), .B1(new_n671_), .B2(new_n398_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT110), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT47), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n704_), .A2(new_n706_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1330gat));
  INV_X1    g510(.A(G50gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n671_), .A2(new_n712_), .A3(new_n555_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n680_), .A2(new_n714_), .A3(new_n555_), .A4(new_n681_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(G50gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n680_), .A2(new_n555_), .A3(new_n681_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT111), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n716_), .A2(KEYINPUT112), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT112), .B1(new_n716_), .B2(new_n718_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n713_), .B1(new_n719_), .B2(new_n720_), .ZN(G1331gat));
  AOI21_X1  g520(.A(new_n296_), .B1(new_n557_), .B2(new_n576_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n262_), .A2(new_n265_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n642_), .A4(new_n625_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n441_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n627_), .A2(new_n723_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT113), .Z(new_n727_));
  INV_X1    g526(.A(new_n296_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n641_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n722_), .A2(KEYINPUT114), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n727_), .A2(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n441_), .A2(G57gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n725_), .B1(new_n734_), .B2(new_n735_), .ZN(G1332gat));
  OAI21_X1  g535(.A(G64gat), .B1(new_n724_), .B2(new_n647_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT48), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n647_), .A2(G64gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n734_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(G1333gat));
  OAI21_X1  g541(.A(G71gat), .B1(new_n724_), .B2(new_n655_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT49), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n655_), .A2(G71gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n734_), .B2(new_n745_), .ZN(G1334gat));
  OAI21_X1  g545(.A(G78gat), .B1(new_n724_), .B2(new_n490_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT50), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n490_), .A2(G78gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n734_), .B2(new_n749_), .ZN(G1335gat));
  INV_X1    g549(.A(new_n723_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(new_n669_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n733_), .A2(KEYINPUT116), .A3(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n440_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT117), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n759_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n674_), .A2(new_n677_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n751_), .A2(new_n296_), .A3(new_n625_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT118), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n441_), .A2(new_n215_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n760_), .A2(new_n761_), .B1(new_n765_), .B2(new_n766_), .ZN(G1336gat));
  AOI21_X1  g566(.A(G92gat), .B1(new_n757_), .B2(new_n554_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT119), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n769_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n647_), .A2(new_n216_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(new_n770_), .A2(new_n771_), .B1(new_n765_), .B2(new_n772_), .ZN(G1337gat));
  AND2_X1   g572(.A1(new_n398_), .A2(new_n210_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n762_), .A2(new_n398_), .A3(new_n763_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n757_), .A2(new_n774_), .B1(G99gat), .B2(new_n775_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g576(.A1(new_n762_), .A2(new_n555_), .A3(new_n763_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G106gat), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT52), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n781_), .A3(G106gat), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n490_), .A2(G106gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n757_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n785_), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT120), .B(new_n787_), .C1(new_n753_), .C2(new_n756_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n783_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n783_), .B(new_n791_), .C1(new_n786_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n283_), .A2(G229gat), .A3(G233gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n293_), .B1(new_n286_), .B2(new_n284_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n288_), .A2(new_n293_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n264_), .B2(new_n259_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n249_), .B2(new_n203_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n249_), .A2(new_n203_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n249_), .A2(new_n799_), .A3(new_n203_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n245_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT56), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n245_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n805_), .A2(new_n296_), .A3(new_n256_), .A4(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n798_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT121), .B(new_n794_), .C1(new_n809_), .C2(new_n667_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n667_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT57), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n805_), .A2(new_n256_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n797_), .A3(new_n807_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n814_), .A2(KEYINPUT58), .A3(new_n797_), .A4(new_n807_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n676_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n813_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n668_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n296_), .B(new_n668_), .C1(new_n606_), .C2(new_n608_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n265_), .A3(new_n262_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n821_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n828_));
  OR3_X1    g627(.A1(new_n640_), .A2(new_n828_), .A3(new_n441_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n640_), .B2(new_n441_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n296_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT59), .B1(new_n827_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n832_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n827_), .B(new_n831_), .C1(new_n836_), .C2(KEYINPUT59), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n728_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n835_), .B1(new_n840_), .B2(new_n834_), .ZN(G1340gat));
  INV_X1    g640(.A(G120gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n751_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n833_), .B(new_n843_), .C1(KEYINPUT60), .C2(new_n842_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n751_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n842_), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n833_), .A2(new_n847_), .A3(new_n625_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n668_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1342gat));
  NAND2_X1  g649(.A1(new_n676_), .A2(G134gat), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n825_), .B1(new_n820_), .B2(new_n668_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n831_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n854_), .A2(new_n642_), .A3(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n853_), .B1(new_n856_), .B2(G134gat), .ZN(new_n857_));
  INV_X1    g656(.A(G134gat), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT124), .B(new_n858_), .C1(new_n832_), .C2(new_n642_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n852_), .A2(new_n860_), .ZN(G1343gat));
  NAND4_X1  g660(.A1(new_n655_), .A2(new_n440_), .A3(new_n647_), .A4(new_n555_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n854_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n296_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT125), .B(G141gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1344gat));
  NAND2_X1  g665(.A1(new_n863_), .A2(new_n723_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n625_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  INV_X1    g670(.A(new_n863_), .ZN(new_n872_));
  OR3_X1    g671(.A1(new_n872_), .A2(G162gat), .A3(new_n642_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G162gat), .B1(new_n872_), .B2(new_n609_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1347gat));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n854_), .A2(new_n647_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n655_), .A2(new_n440_), .A3(new_n555_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n877_), .A2(new_n296_), .A3(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n876_), .B1(new_n879_), .B2(new_n304_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n878_), .ZN(new_n881_));
  OAI211_X1 g680(.A(KEYINPUT62), .B(G169gat), .C1(new_n881_), .C2(new_n728_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n879_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n882_), .A3(new_n883_), .ZN(G1348gat));
  NAND3_X1  g683(.A1(new_n877_), .A2(new_n723_), .A3(new_n878_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g685(.A1(new_n877_), .A2(new_n625_), .A3(new_n878_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n512_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n312_), .B2(new_n887_), .ZN(G1350gat));
  OAI21_X1  g688(.A(G190gat), .B1(new_n881_), .B2(new_n609_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n667_), .A2(new_n511_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n881_), .B2(new_n891_), .ZN(G1351gat));
  NOR3_X1   g691(.A1(new_n398_), .A2(new_n440_), .A3(new_n490_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n877_), .A2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n448_), .B1(new_n894_), .B2(new_n728_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n877_), .A2(G197gat), .A3(new_n296_), .A4(new_n893_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n827_), .A2(new_n554_), .A3(new_n893_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n899_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n296_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n895_), .A2(new_n898_), .A3(new_n900_), .ZN(G1352gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n723_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n894_), .B2(new_n668_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT63), .B(G211gat), .Z(new_n906_));
  NAND4_X1  g705(.A1(new_n877_), .A2(new_n625_), .A3(new_n893_), .A4(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT127), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n899_), .A2(new_n909_), .A3(new_n625_), .A4(new_n906_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n905_), .A2(new_n908_), .A3(new_n910_), .ZN(G1354gat));
  OAI21_X1  g710(.A(G218gat), .B1(new_n894_), .B2(new_n609_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n899_), .A2(new_n455_), .A3(new_n667_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1355gat));
endmodule


