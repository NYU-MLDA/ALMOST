//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_;
  INV_X1    g000(.A(G183gat), .ZN(new_n202_));
  INV_X1    g001(.A(G190gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT23), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT87), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(KEYINPUT87), .A3(new_n210_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n208_), .A2(new_n213_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT86), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n206_), .A2(new_n217_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n205_), .A2(KEYINPUT86), .A3(G183gat), .A4(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n204_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT85), .B1(new_n203_), .B2(KEYINPUT26), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT85), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(G183gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n202_), .A2(KEYINPUT84), .A3(KEYINPUT25), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n203_), .A2(KEYINPUT26), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(G183gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n226_), .A2(new_n231_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT24), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(G169gat), .B2(G176gat), .ZN(new_n237_));
  OR2_X1    g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n235_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n221_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n216_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n241_), .B(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  XOR2_X1   g045(.A(G127gat), .B(G134gat), .Z(new_n247_));
  XOR2_X1   g046(.A(G113gat), .B(G120gat), .Z(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(G15gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT30), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n249_), .B(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n246_), .B(new_n254_), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT89), .ZN(new_n256_));
  INV_X1    g055(.A(G218gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G211gat), .ZN(new_n258_));
  INV_X1    g057(.A(G211gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G218gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n260_), .A3(KEYINPUT94), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT94), .B1(new_n258_), .B2(new_n260_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT95), .ZN(new_n265_));
  INV_X1    g064(.A(G204gat), .ZN(new_n266_));
  INV_X1    g065(.A(G197gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT93), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT93), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G197gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n266_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G197gat), .A2(G204gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n265_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n272_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT93), .B(G197gat), .ZN(new_n275_));
  OAI211_X1 g074(.A(KEYINPUT95), .B(new_n274_), .C1(new_n275_), .C2(new_n266_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n264_), .A2(new_n273_), .A3(KEYINPUT21), .A4(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n258_), .A2(new_n260_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT94), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n261_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n275_), .A2(new_n266_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n278_), .B1(G197gat), .B2(G204gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n279_), .A2(new_n283_), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n277_), .A2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT20), .B1(new_n288_), .B2(new_n241_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n224_), .A2(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n202_), .A2(KEYINPUT25), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n239_), .A2(new_n207_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT98), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT99), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n214_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT99), .A2(G169gat), .A3(G176gat), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n209_), .A2(new_n210_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n205_), .B1(G183gat), .B2(G190gat), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n298_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT98), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n239_), .A2(new_n303_), .A3(new_n207_), .A4(new_n292_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n294_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n288_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT100), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT100), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n288_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n289_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT19), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n277_), .A2(new_n287_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(new_n302_), .A3(new_n293_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT20), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n288_), .B2(new_n241_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n312_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G8gat), .B(G36gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G64gat), .B(G92gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT106), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n318_), .B(new_n313_), .C1(new_n288_), .C2(new_n305_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n326_), .B(new_n329_), .C1(new_n310_), .C2(new_n313_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(KEYINPUT27), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT107), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n329_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n326_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n330_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT27), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n332_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  AOI211_X1 g137(.A(KEYINPUT107), .B(KEYINPUT27), .C1(new_n335_), .C2(new_n330_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n331_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G228gat), .A2(G233gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  INV_X1    g142(.A(G155gat), .ZN(new_n344_));
  INV_X1    g143(.A(G162gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT90), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT90), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(G155gat), .A3(G162gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n343_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n349_), .A2(KEYINPUT92), .ZN(new_n350_));
  OR3_X1    g149(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .A4(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n349_), .B2(KEYINPUT92), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n350_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT91), .ZN(new_n360_));
  INV_X1    g159(.A(G141gat), .ZN(new_n361_));
  INV_X1    g160(.A(G148gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n352_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n346_), .A2(new_n348_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n343_), .B1(new_n365_), .B2(KEYINPUT1), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n346_), .A2(new_n367_), .A3(new_n348_), .ZN(new_n368_));
  AOI211_X1 g167(.A(new_n360_), .B(new_n364_), .C1(new_n366_), .C2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(KEYINPUT1), .ZN(new_n370_));
  INV_X1    g169(.A(new_n343_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n364_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT91), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n359_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT29), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n342_), .B1(new_n376_), .B2(new_n288_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n342_), .ZN(new_n378_));
  AOI211_X1 g177(.A(new_n315_), .B(new_n378_), .C1(new_n375_), .C2(KEYINPUT29), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n341_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n350_), .A2(new_n358_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n346_), .A2(new_n367_), .A3(new_n348_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n367_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n343_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n360_), .B1(new_n384_), .B2(new_n364_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n372_), .A2(KEYINPUT91), .A3(new_n373_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n381_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n288_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n378_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n376_), .A2(new_n288_), .A3(new_n342_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n341_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT96), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n380_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G22gat), .B(G50gat), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n388_), .B(new_n359_), .C1(new_n369_), .C2(new_n374_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT28), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n385_), .A2(new_n386_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n388_), .A4(new_n359_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n396_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n398_), .A2(new_n401_), .A3(new_n396_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT96), .B(new_n341_), .C1(new_n377_), .C2(new_n379_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n398_), .A2(new_n401_), .A3(new_n396_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(new_n402_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT97), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n390_), .A2(new_n391_), .A3(new_n410_), .A4(new_n392_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n411_), .A3(new_n380_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n393_), .A2(KEYINPUT97), .ZN(new_n413_));
  OAI22_X1  g212(.A1(new_n395_), .A2(new_n407_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n375_), .A2(new_n249_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n249_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n399_), .A2(new_n416_), .A3(new_n359_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n417_), .A3(KEYINPUT4), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n375_), .A2(new_n421_), .A3(new_n249_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n418_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n415_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT103), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT103), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n415_), .A2(new_n417_), .A3(new_n426_), .A4(new_n419_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G1gat), .B(G29gat), .Z(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n423_), .A2(new_n425_), .A3(new_n435_), .A4(new_n427_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n414_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n340_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(KEYINPUT104), .A2(KEYINPUT33), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n440_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n415_), .A2(new_n417_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n433_), .B1(new_n443_), .B2(new_n419_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT105), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n418_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT105), .B(new_n433_), .C1(new_n443_), .C2(new_n419_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n335_), .A2(new_n330_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n441_), .A2(new_n442_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n434_), .A2(new_n436_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n321_), .A2(KEYINPUT32), .A3(new_n326_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n454_), .B(new_n329_), .C1(new_n310_), .C2(new_n313_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n414_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n256_), .B1(new_n439_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n340_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n414_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n459_), .A2(new_n255_), .A3(new_n437_), .A4(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT13), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT72), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT70), .ZN(new_n465_));
  XOR2_X1   g264(.A(G85gat), .B(G92gat), .Z(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(G99gat), .B2(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(KEYINPUT6), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT69), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(KEYINPUT6), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n467_), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT69), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT68), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n481_));
  INV_X1    g280(.A(G99gat), .ZN(new_n482_));
  INV_X1    g281(.A(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n477_), .B1(new_n481_), .B2(KEYINPUT68), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n480_), .A2(new_n481_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n466_), .B1(new_n476_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n472_), .A2(new_n473_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT66), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT66), .B1(new_n472_), .B2(new_n473_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT7), .B1(new_n478_), .B2(new_n479_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT67), .B1(new_n479_), .B2(KEYINPUT7), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(new_n484_), .ZN(new_n495_));
  OAI22_X1  g294(.A1(new_n491_), .A2(new_n492_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n466_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n488_), .A2(KEYINPUT8), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n483_), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT64), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n489_), .B(new_n490_), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT65), .B(G85gat), .Z(new_n506_));
  INV_X1    g305(.A(G92gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(KEYINPUT9), .ZN(new_n508_));
  AOI22_X1  g307(.A1(KEYINPUT9), .A2(new_n466_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n465_), .B1(new_n500_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G57gat), .B(G64gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT11), .Z(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT71), .B(G71gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(G78gat), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(KEYINPUT11), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n471_), .B(new_n475_), .C1(new_n493_), .C2(new_n495_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n497_), .B1(new_n521_), .B2(new_n466_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT68), .B1(new_n484_), .B2(new_n477_), .ZN(new_n523_));
  OAI22_X1  g322(.A1(new_n523_), .A2(KEYINPUT7), .B1(new_n484_), .B2(new_n494_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n498_), .B1(new_n505_), .B2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(KEYINPUT70), .B(new_n510_), .C1(new_n522_), .C2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n512_), .A2(new_n520_), .A3(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n510_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n517_), .A2(new_n519_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(KEYINPUT12), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n520_), .B1(new_n512_), .B2(new_n526_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n527_), .B(new_n530_), .C1(new_n531_), .C2(KEYINPUT12), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G230gat), .A2(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n464_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n526_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n496_), .A2(new_n499_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n466_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n474_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n541_), .B2(new_n524_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n537_), .B1(new_n542_), .B2(new_n497_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT70), .B1(new_n543_), .B2(new_n510_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n529_), .B1(new_n536_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n527_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n534_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n527_), .A2(new_n530_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n548_), .A2(new_n550_), .A3(KEYINPUT72), .A4(new_n533_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n535_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G120gat), .B(G148gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT5), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G176gat), .B(G204gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n535_), .A2(new_n551_), .A3(new_n547_), .A4(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(KEYINPUT73), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT73), .B1(new_n557_), .B2(new_n559_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n463_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n557_), .A2(new_n559_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT73), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(KEYINPUT13), .A3(new_n560_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G29gat), .B(G36gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G43gat), .B(G50gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT15), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573_));
  INV_X1    g372(.A(G1gat), .ZN(new_n574_));
  INV_X1    g373(.A(G8gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G1gat), .B(G8gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n572_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n571_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n579_), .B(new_n571_), .Z(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(G229gat), .A3(G233gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT81), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G169gat), .B(G197gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT82), .ZN(new_n594_));
  INV_X1    g393(.A(new_n592_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n585_), .A2(new_n587_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n588_), .A2(KEYINPUT82), .A3(new_n592_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT83), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT83), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n462_), .A2(new_n568_), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT35), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n512_), .A2(new_n571_), .A3(new_n526_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT74), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT74), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n512_), .A2(new_n619_), .A3(new_n571_), .A4(new_n526_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n528_), .A2(new_n572_), .B1(new_n614_), .B2(new_n613_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n616_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n615_), .B(new_n624_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n610_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT75), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  OAI221_X1 g430(.A(new_n627_), .B1(new_n629_), .B2(new_n610_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT76), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT77), .B1(new_n631_), .B2(new_n632_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n635_), .B(KEYINPUT37), .C1(new_n634_), .C2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT77), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n634_), .B1(new_n633_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n579_), .B(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n520_), .B(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G127gat), .B(G155gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G183gat), .B(G211gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT17), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n645_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT79), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n650_), .A2(KEYINPUT17), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n645_), .A2(new_n651_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT80), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT80), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n642_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n606_), .A2(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n661_), .A2(new_n574_), .A3(new_n452_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT38), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT108), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n458_), .A2(new_n461_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n633_), .B(KEYINPUT109), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n656_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n568_), .A2(new_n599_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n670_), .B2(new_n437_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n664_), .B(new_n671_), .C1(KEYINPUT38), .C2(new_n662_), .ZN(G1324gat));
  NAND3_X1  g471(.A1(new_n661_), .A2(new_n575_), .A3(new_n340_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n340_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n676_), .B2(G8gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(G8gat), .B1(new_n670_), .B2(new_n459_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(KEYINPUT39), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n673_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT111), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT111), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n673_), .C1(new_n677_), .C2(new_n679_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n681_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  INV_X1    g486(.A(new_n256_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n251_), .B1(new_n675_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT41), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n661_), .A2(new_n251_), .A3(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT112), .ZN(G1326gat));
  XNOR2_X1  g492(.A(new_n414_), .B(KEYINPUT113), .ZN(new_n694_));
  OAI21_X1  g493(.A(G22gat), .B1(new_n670_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT42), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n694_), .A2(G22gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT114), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n661_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1327gat));
  INV_X1    g499(.A(new_n659_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n633_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n606_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n452_), .ZN(new_n706_));
  AOI221_X4 g505(.A(KEYINPUT43), .B1(new_n458_), .B2(new_n461_), .C1(new_n637_), .C2(new_n641_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n642_), .B2(new_n665_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n669_), .A2(new_n659_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n452_), .A2(G29gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n706_), .B1(new_n715_), .B2(new_n716_), .ZN(G1328gat));
  NAND3_X1  g516(.A1(new_n713_), .A2(new_n340_), .A3(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G36gat), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n704_), .A2(G36gat), .A3(new_n459_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT45), .Z(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n721_), .A3(KEYINPUT46), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1329gat));
  NAND4_X1  g525(.A1(new_n713_), .A2(G43gat), .A3(new_n255_), .A4(new_n714_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n704_), .A2(new_n256_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(G43gat), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g529(.A(new_n694_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G50gat), .B1(new_n705_), .B2(new_n731_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n414_), .A2(G50gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n715_), .B2(new_n733_), .ZN(G1331gat));
  NOR2_X1   g533(.A1(new_n659_), .A2(new_n604_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n568_), .A2(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n667_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G57gat), .B1(new_n738_), .B2(new_n437_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n568_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n462_), .A2(new_n740_), .A3(new_n600_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n660_), .ZN(new_n742_));
  INV_X1    g541(.A(G57gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n452_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n739_), .A2(new_n744_), .ZN(G1332gat));
  INV_X1    g544(.A(G64gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n737_), .B2(new_n340_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT48), .Z(new_n748_));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n746_), .A3(new_n340_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1333gat));
  INV_X1    g549(.A(G71gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n737_), .B2(new_n688_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT49), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n742_), .A2(new_n751_), .A3(new_n688_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1334gat));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n737_), .B2(new_n731_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n742_), .A2(new_n756_), .A3(new_n731_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1335gat));
  NAND2_X1  g560(.A1(new_n741_), .A2(new_n703_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G85gat), .B1(new_n763_), .B2(new_n452_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n636_), .A2(new_n634_), .A3(KEYINPUT37), .ZN(new_n765_));
  INV_X1    g564(.A(new_n639_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n640_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n768_), .B2(new_n462_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n642_), .A2(new_n708_), .A3(new_n665_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n561_), .A2(new_n562_), .A3(new_n463_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT13), .B1(new_n566_), .B2(new_n560_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n659_), .B(new_n599_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n568_), .A2(KEYINPUT116), .A3(new_n659_), .A4(new_n599_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n769_), .A2(new_n770_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n452_), .A2(new_n506_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n764_), .B1(new_n777_), .B2(new_n778_), .ZN(G1336gat));
  AOI21_X1  g578(.A(G92gat), .B1(new_n763_), .B2(new_n340_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n340_), .A2(G92gat), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT117), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n777_), .B2(new_n782_), .ZN(G1337gat));
  AND4_X1   g582(.A1(new_n501_), .A2(new_n763_), .A3(new_n502_), .A4(new_n255_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n482_), .B1(new_n777_), .B2(new_n688_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT51), .Z(G1338gat));
  NAND2_X1  g586(.A1(new_n775_), .A2(new_n776_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n788_), .B(new_n414_), .C1(new_n709_), .C2(new_n707_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n790_));
  OAI21_X1  g589(.A(G106gat), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT118), .B1(new_n777_), .B2(new_n414_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT52), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n790_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n777_), .A2(KEYINPUT118), .A3(new_n414_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .A4(G106gat), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n793_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n763_), .A2(new_n483_), .A3(new_n414_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n798_), .A2(new_n802_), .A3(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1339gat));
  AOI21_X1  g603(.A(new_n595_), .B1(new_n586_), .B2(new_n584_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n583_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n584_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n596_), .A2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n559_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n548_), .A2(new_n550_), .A3(KEYINPUT55), .A4(new_n533_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT121), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n810_), .A2(new_n811_), .B1(new_n534_), .B2(new_n532_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n535_), .A2(new_n814_), .A3(new_n551_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n816_), .A2(KEYINPUT56), .A3(new_n556_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT56), .B1(new_n816_), .B2(new_n556_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n809_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n820_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n642_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n600_), .A2(new_n559_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n600_), .A2(KEYINPUT120), .A3(new_n559_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n827_), .B(new_n828_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n808_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n824_), .B1(new_n831_), .B2(new_n702_), .ZN(new_n832_));
  AOI211_X1 g631(.A(KEYINPUT57), .B(new_n633_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n823_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n659_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n768_), .A2(new_n740_), .A3(new_n735_), .A4(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n836_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n735_), .A2(new_n567_), .A3(new_n563_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n642_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n835_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  AND4_X1   g643(.A1(new_n255_), .A2(new_n459_), .A3(new_n452_), .A4(new_n460_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n834_), .A2(new_n656_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n842_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n845_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n846_), .B1(new_n850_), .B2(new_n844_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n605_), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n849_), .A2(G113gat), .A3(new_n599_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n851_), .B2(new_n740_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n740_), .A2(KEYINPUT60), .ZN(new_n856_));
  MUX2_X1   g655(.A(new_n856_), .B(KEYINPUT60), .S(G120gat), .Z(new_n857_));
  NAND2_X1  g656(.A1(new_n850_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(G1341gat));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n849_), .B2(new_n659_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n849_), .A2(KEYINPUT59), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT123), .B(G127gat), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n864_), .A2(new_n668_), .A3(new_n846_), .A4(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n863_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n861_), .A2(new_n862_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1342gat));
  OAI21_X1  g668(.A(G134gat), .B1(new_n851_), .B2(new_n768_), .ZN(new_n870_));
  OR3_X1    g669(.A1(new_n849_), .A2(G134gat), .A3(new_n666_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1343gat));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n841_), .B1(new_n834_), .B2(new_n656_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n688_), .A2(new_n460_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n459_), .A2(new_n452_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n873_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n874_), .A2(KEYINPUT124), .A3(new_n876_), .A4(new_n878_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n600_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G141gat), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n361_), .B(new_n600_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1344gat));
  OAI21_X1  g684(.A(new_n568_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G148gat), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n362_), .B(new_n568_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1345gat));
  OAI21_X1  g688(.A(new_n701_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n891_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n701_), .B(new_n893_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1346gat));
  INV_X1    g694(.A(new_n666_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n345_), .B(new_n896_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n881_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n848_), .A2(new_n875_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT124), .B1(new_n899_), .B2(new_n878_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n768_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n897_), .B1(new_n901_), .B2(new_n345_), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n459_), .A2(new_n452_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n256_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n731_), .A2(new_n599_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n843_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G169gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT125), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n907_), .A2(new_n910_), .A3(G169gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n909_), .A2(KEYINPUT62), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n908_), .A2(KEYINPUT125), .A3(new_n913_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n843_), .A2(new_n209_), .A3(new_n905_), .A4(new_n906_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n912_), .A2(new_n914_), .A3(new_n915_), .ZN(G1348gat));
  AND3_X1   g715(.A1(new_n843_), .A2(new_n694_), .A3(new_n905_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G176gat), .B1(new_n917_), .B2(new_n568_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n874_), .A2(new_n414_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n905_), .A2(G176gat), .A3(new_n568_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1349gat));
  NAND3_X1  g720(.A1(new_n919_), .A2(new_n701_), .A3(new_n905_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n656_), .B1(new_n291_), .B2(new_n233_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n922_), .A2(new_n202_), .B1(new_n917_), .B2(new_n923_), .ZN(G1350gat));
  AND3_X1   g723(.A1(new_n896_), .A2(new_n290_), .A3(new_n232_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n917_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n843_), .A2(new_n694_), .A3(new_n905_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G190gat), .B1(new_n927_), .B2(new_n768_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT126), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n926_), .A2(new_n928_), .A3(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1351gat));
  NOR2_X1   g732(.A1(new_n899_), .A2(new_n904_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n600_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT127), .B(G197gat), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1352gat));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n568_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g738(.A1(new_n899_), .A2(new_n656_), .A3(new_n904_), .ZN(new_n940_));
  OR2_X1    g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  XOR2_X1   g741(.A(KEYINPUT63), .B(G211gat), .Z(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n940_), .B2(new_n943_), .ZN(G1354gat));
  NAND3_X1  g743(.A1(new_n934_), .A2(new_n257_), .A3(new_n896_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n899_), .A2(new_n768_), .A3(new_n904_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(new_n257_), .ZN(G1355gat));
endmodule


