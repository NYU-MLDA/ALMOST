//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n203_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT3), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(G141gat), .B2(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(KEYINPUT76), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n208_), .A2(KEYINPUT76), .A3(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n202_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n214_), .A2(new_n216_), .A3(KEYINPUT77), .A4(new_n218_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n210_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G134gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G127gat), .ZN(new_n225_));
  INV_X1    g024(.A(G127gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G134gat), .ZN(new_n227_));
  AND3_X1   g026(.A1(new_n225_), .A2(new_n227_), .A3(KEYINPUT74), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT74), .B1(new_n225_), .B2(new_n227_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G113gat), .B(G120gat), .Z(new_n230_));
  NOR3_X1   g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT74), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n226_), .A2(G134gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n224_), .A2(G127gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n225_), .A2(new_n227_), .A3(KEYINPUT74), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n232_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT89), .B1(new_n231_), .B2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n230_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n237_), .A3(new_n232_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT89), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n223_), .A2(KEYINPUT90), .A3(new_n239_), .A4(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n210_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n219_), .A2(new_n220_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n202_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n222_), .ZN(new_n248_));
  AND4_X1   g047(.A1(new_n245_), .A2(new_n239_), .A3(new_n248_), .A4(new_n243_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT90), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n231_), .A2(new_n238_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n223_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n244_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G1gat), .B(G29gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G57gat), .B(G85gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n248_), .A2(new_n245_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n251_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n223_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n250_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n262_), .B1(new_n267_), .B2(new_n244_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n254_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n255_), .B(new_n261_), .C1(new_n268_), .C2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT33), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n253_), .A2(KEYINPUT4), .ZN(new_n274_));
  INV_X1    g073(.A(new_n271_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT33), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n261_), .A4(new_n255_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n253_), .A2(new_n270_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n260_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n269_), .A2(new_n254_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n253_), .B2(KEYINPUT4), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT92), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n261_), .B1(new_n253_), .B2(new_n270_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT92), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n284_), .B(new_n285_), .C1(new_n268_), .C2(new_n281_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n273_), .A2(new_n278_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G8gat), .B(G36gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT18), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G64gat), .B(G92gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT19), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT20), .ZN(new_n296_));
  OR2_X1    g095(.A1(KEYINPUT80), .A2(G197gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(KEYINPUT80), .A2(G197gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(G204gat), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT82), .ZN(new_n300_));
  AND2_X1   g099(.A1(KEYINPUT81), .A2(G204gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(KEYINPUT81), .A2(G204gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n304_), .A3(G197gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n297_), .A2(new_n306_), .A3(G204gat), .A4(new_n298_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n300_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G211gat), .B(G218gat), .Z(new_n309_));
  AND2_X1   g108(.A1(new_n309_), .A2(KEYINPUT21), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(G204gat), .ZN(new_n313_));
  AND2_X1   g112(.A1(KEYINPUT80), .A2(G197gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(KEYINPUT80), .A2(G197gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G197gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n309_), .B1(new_n319_), .B2(KEYINPUT21), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT83), .B(KEYINPUT21), .Z(new_n321_));
  NAND4_X1  g120(.A1(new_n300_), .A2(new_n305_), .A3(new_n307_), .A4(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT84), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n320_), .A2(new_n322_), .A3(KEYINPUT84), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n312_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT23), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(G183gat), .B2(G190gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(KEYINPUT70), .A2(G169gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(G176gat), .B1(new_n333_), .B2(KEYINPUT22), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT22), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT70), .A3(G169gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n332_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n330_), .B1(new_n338_), .B2(KEYINPUT71), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT24), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT25), .B(G183gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT26), .B(G190gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n348_), .A3(new_n329_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n331_), .A2(KEYINPUT24), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n349_), .B1(new_n344_), .B2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n342_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n296_), .B1(new_n327_), .B2(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n320_), .A2(new_n322_), .A3(KEYINPUT84), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT84), .B1(new_n320_), .B2(new_n322_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n311_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n344_), .B1(new_n351_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n350_), .A2(KEYINPUT87), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n349_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G169gat), .ZN(new_n364_));
  INV_X1    g163(.A(G176gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n332_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n362_), .A2(new_n363_), .B1(new_n330_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n357_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n295_), .B1(new_n354_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT20), .B1(new_n327_), .B2(new_n353_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n295_), .B1(new_n357_), .B2(new_n368_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n292_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n363_), .B1(new_n343_), .B2(new_n350_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n341_), .B2(new_n339_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT20), .B1(new_n357_), .B2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n327_), .A2(new_n367_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n294_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n294_), .B1(new_n327_), .B2(new_n367_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n296_), .B1(new_n357_), .B2(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n291_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n374_), .A2(KEYINPUT88), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n385_), .B(new_n292_), .C1(new_n370_), .C2(new_n373_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n287_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n276_), .A2(new_n255_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n260_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n272_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n291_), .A2(KEYINPUT32), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n367_), .A2(KEYINPUT93), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n330_), .A2(new_n366_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n394_), .B(KEYINPUT93), .C1(new_n361_), .C2(new_n349_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n393_), .A2(new_n357_), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n294_), .B1(new_n397_), .B2(new_n371_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n354_), .A2(new_n295_), .A3(new_n369_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n392_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n379_), .A2(new_n382_), .A3(new_n392_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n391_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n388_), .A2(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT78), .B(KEYINPUT28), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n248_), .A2(new_n407_), .A3(new_n245_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G22gat), .B(G50gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n409_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n223_), .B2(new_n407_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n406_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n409_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n223_), .A2(new_n407_), .A3(new_n411_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n405_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(KEYINPUT79), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(KEYINPUT79), .A2(G233gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(G228gat), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n223_), .A2(new_n407_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n425_), .B1(new_n327_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n263_), .A2(KEYINPUT29), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n357_), .A2(new_n428_), .A3(new_n424_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n420_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n418_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT86), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n327_), .A2(new_n426_), .A3(new_n425_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n424_), .B1(new_n357_), .B2(new_n428_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n419_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT85), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n418_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n434_), .A2(new_n435_), .A3(new_n419_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n430_), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n433_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(new_n433_), .B2(new_n439_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n441_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n438_), .B1(new_n437_), .B2(new_n418_), .ZN(new_n446_));
  AOI211_X1 g245(.A(KEYINPUT86), .B(new_n417_), .C1(new_n436_), .C2(KEYINPUT85), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n433_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n391_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT27), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n384_), .A2(new_n451_), .A3(new_n386_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n398_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n399_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n292_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(KEYINPUT27), .A3(new_n383_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n404_), .A2(new_n444_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n376_), .B(KEYINPUT30), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT73), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n460_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G227gat), .A2(G233gat), .ZN(new_n463_));
  INV_X1    g262(.A(G15gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G71gat), .ZN(new_n466_));
  INV_X1    g265(.A(G99gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(KEYINPUT72), .B(G43gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n461_), .A2(new_n462_), .A3(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n251_), .B(KEYINPUT31), .Z(new_n472_));
  INV_X1    g271(.A(KEYINPUT75), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n471_), .B(new_n474_), .C1(new_n462_), .C2(new_n470_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n472_), .A2(new_n473_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT94), .B1(new_n458_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n448_), .A2(new_n449_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n452_), .A2(new_n456_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n391_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n287_), .A2(new_n387_), .B1(new_n391_), .B2(new_n402_), .ZN(new_n485_));
  OAI22_X1  g284(.A1(new_n484_), .A2(new_n480_), .B1(new_n485_), .B2(new_n479_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n487_));
  INV_X1    g286(.A(new_n477_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n478_), .A2(new_n483_), .A3(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G29gat), .B(G36gat), .Z(new_n491_));
  XOR2_X1   g290(.A(G43gat), .B(G50gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT15), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495_));
  INV_X1    g294(.A(G1gat), .ZN(new_n496_));
  INV_X1    g295(.A(G8gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT14), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G1gat), .B(G8gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n494_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n493_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n501_), .B(new_n493_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n508_), .B2(new_n505_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G169gat), .B(G197gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n509_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT69), .Z(new_n514_));
  AND2_X1   g313(.A1(new_n490_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G85gat), .B(G92gat), .Z(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(KEYINPUT9), .B2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT10), .B(G99gat), .Z(new_n521_));
  INV_X1    g320(.A(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT64), .B(G92gat), .Z(new_n524_));
  INV_X1    g323(.A(KEYINPUT9), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(G85gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n520_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT7), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n519_), .B1(new_n530_), .B2(new_n518_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n531_), .A2(KEYINPUT8), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(KEYINPUT8), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n527_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n537_));
  XOR2_X1   g336(.A(G71gat), .B(G78gat), .Z(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n537_), .A2(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n534_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n541_), .B(new_n527_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(KEYINPUT12), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT12), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n534_), .A2(new_n546_), .A3(new_n542_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT65), .ZN(new_n551_));
  INV_X1    g350(.A(new_n549_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT65), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n543_), .A2(new_n544_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n551_), .B(new_n555_), .C1(new_n549_), .C2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT5), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n557_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT13), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT66), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(KEYINPUT66), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n541_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT68), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n501_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G127gat), .B(G155gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT16), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n575_), .A2(new_n576_), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n571_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n571_), .A2(new_n577_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n494_), .A2(new_n534_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  INV_X1    g383(.A(new_n493_), .ZN(new_n585_));
  OAI221_X1 g384(.A(new_n582_), .B1(KEYINPUT35), .B2(new_n584_), .C1(new_n585_), .C2(new_n534_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT67), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n586_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(KEYINPUT36), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(KEYINPUT36), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n589_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  AND4_X1   g397(.A1(new_n515_), .A2(new_n567_), .A3(new_n581_), .A4(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n496_), .A3(new_n391_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT95), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n596_), .B(KEYINPUT96), .Z(new_n605_));
  AND2_X1   g404(.A1(new_n490_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n606_), .A2(new_n567_), .A3(new_n514_), .A4(new_n581_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT97), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT97), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n482_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n603_), .B(new_n604_), .C1(new_n496_), .C2(new_n610_), .ZN(G1324gat));
  OAI21_X1  g410(.A(G8gat), .B1(new_n607_), .B2(new_n457_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT39), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n599_), .A2(new_n497_), .A3(new_n480_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n608_), .A2(new_n609_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n477_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n619_), .B2(G15gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI211_X1 g420(.A(KEYINPUT98), .B(new_n464_), .C1(new_n618_), .C2(new_n477_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n623_), .A3(KEYINPUT41), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n599_), .A2(new_n464_), .A3(new_n477_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n626_), .A3(new_n627_), .ZN(G1326gat));
  INV_X1    g427(.A(G22gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n618_), .B2(new_n479_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT99), .B(KEYINPUT42), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n599_), .A2(new_n629_), .A3(new_n479_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1327gat));
  INV_X1    g433(.A(new_n581_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(new_n596_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n515_), .A2(new_n567_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n515_), .A2(new_n567_), .A3(KEYINPUT102), .A4(new_n636_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(G29gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n391_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n514_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n566_), .A2(new_n644_), .A3(new_n581_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n598_), .B1(new_n490_), .B2(KEYINPUT100), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n478_), .A2(new_n648_), .A3(new_n483_), .A4(new_n489_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n646_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n598_), .A2(KEYINPUT43), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n489_), .A2(new_n483_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n487_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT101), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n490_), .A2(new_n656_), .A3(new_n651_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n645_), .B1(new_n650_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT44), .B(new_n645_), .C1(new_n650_), .C2(new_n658_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n661_), .A2(new_n391_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n643_), .B1(new_n663_), .B2(new_n642_), .ZN(G1328gat));
  NOR2_X1   g463(.A1(new_n457_), .A2(G36gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n639_), .A2(new_n640_), .A3(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT45), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n661_), .A2(new_n480_), .A3(new_n662_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(KEYINPUT103), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n661_), .A2(new_n670_), .A3(new_n480_), .A4(new_n662_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G36gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n667_), .B1(new_n669_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n667_), .B(KEYINPUT46), .C1(new_n669_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1329gat));
  NAND3_X1  g476(.A1(new_n639_), .A2(new_n477_), .A3(new_n640_), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT104), .B(G43gat), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT105), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n661_), .A2(G43gat), .A3(new_n477_), .A4(new_n662_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT47), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(new_n685_), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1330gat));
  AND4_X1   g486(.A1(G50gat), .A2(new_n661_), .A3(new_n479_), .A4(new_n662_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G50gat), .B1(new_n641_), .B2(new_n479_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1331gat));
  AND2_X1   g489(.A1(new_n490_), .A2(new_n644_), .ZN(new_n691_));
  AND4_X1   g490(.A1(new_n566_), .A2(new_n691_), .A3(new_n581_), .A4(new_n598_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G57gat), .B1(new_n692_), .B2(new_n391_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT106), .Z(new_n694_));
  NAND4_X1  g493(.A1(new_n606_), .A2(new_n644_), .A3(new_n566_), .A4(new_n581_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT107), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT108), .B(G57gat), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n482_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n694_), .B1(new_n696_), .B2(new_n698_), .ZN(G1332gat));
  NOR2_X1   g498(.A1(new_n457_), .A2(G64gat), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT109), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n692_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n695_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n695_), .A2(new_n703_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n480_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(G64gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n706_), .B2(G64gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n702_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT110), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n712_), .B(new_n702_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1333gat));
  INV_X1    g513(.A(G71gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n696_), .B2(new_n477_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT49), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n692_), .A2(new_n715_), .A3(new_n477_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1334gat));
  INV_X1    g518(.A(G78gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n696_), .B2(new_n479_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n692_), .A2(new_n720_), .A3(new_n479_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1335gat));
  OR2_X1    g524(.A1(new_n650_), .A2(new_n658_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n567_), .A2(new_n514_), .A3(new_n581_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G85gat), .B1(new_n728_), .B2(new_n482_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n691_), .A2(new_n566_), .A3(new_n636_), .ZN(new_n730_));
  INV_X1    g529(.A(G85gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n391_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n729_), .A2(new_n732_), .ZN(G1336gat));
  AOI21_X1  g532(.A(G92gat), .B1(new_n730_), .B2(new_n480_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT112), .Z(new_n735_));
  INV_X1    g534(.A(new_n728_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n480_), .A2(new_n524_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(G1337gat));
  NAND3_X1  g537(.A1(new_n730_), .A2(new_n477_), .A3(new_n521_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT113), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(new_n477_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G99gat), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(G1338gat));
  OAI21_X1  g543(.A(G106gat), .B1(new_n728_), .B2(new_n444_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(KEYINPUT52), .B(G106gat), .C1(new_n728_), .C2(new_n444_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n730_), .A2(new_n522_), .A3(new_n479_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT115), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(new_n748_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT53), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n747_), .A2(new_n753_), .A3(new_n748_), .A4(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1339gat));
  NAND4_X1  g554(.A1(new_n563_), .A2(new_n598_), .A3(new_n644_), .A4(new_n581_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT54), .Z(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n557_), .A2(new_n561_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n551_), .A2(new_n761_), .A3(new_n555_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n545_), .A2(KEYINPUT116), .A3(new_n552_), .A4(new_n547_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n764_), .A2(new_n765_), .B1(KEYINPUT55), .B2(new_n553_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n762_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n762_), .A2(new_n766_), .A3(KEYINPUT117), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n561_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n762_), .A2(new_n766_), .A3(KEYINPUT117), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT117), .B1(new_n762_), .B2(new_n766_), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT56), .B(new_n561_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n514_), .B(new_n760_), .C1(new_n772_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n512_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n509_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n512_), .B1(new_n507_), .B2(new_n505_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(KEYINPUT118), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n505_), .B1(new_n501_), .B2(new_n493_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n503_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(KEYINPUT118), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n779_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n562_), .A2(new_n785_), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n758_), .B(new_n596_), .C1(new_n777_), .C2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n760_), .B(new_n785_), .C1(new_n772_), .C2(new_n776_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n561_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n759_), .B1(new_n794_), .B2(new_n775_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n795_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n785_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n598_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n787_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n795_), .A2(new_n514_), .B1(new_n562_), .B2(new_n785_), .ZN(new_n800_));
  OAI211_X1 g599(.A(KEYINPUT119), .B(new_n758_), .C1(new_n800_), .C2(new_n596_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n758_), .B1(new_n800_), .B2(new_n596_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n801_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n757_), .B1(new_n805_), .B2(new_n635_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n481_), .A2(new_n477_), .A3(new_n391_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n514_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n810_));
  INV_X1    g609(.A(new_n757_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n581_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n797_), .A2(new_n798_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n787_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n802_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n635_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(KEYINPUT121), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT122), .B(new_n810_), .C1(new_n814_), .C2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT59), .B1(new_n806_), .B2(new_n807_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(KEYINPUT121), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n812_), .A2(new_n813_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n811_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT122), .B1(new_n825_), .B2(new_n810_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n514_), .A2(G113gat), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT123), .Z(new_n829_));
  AOI21_X1  g628(.A(new_n809_), .B1(new_n827_), .B2(new_n829_), .ZN(G1340gat));
  INV_X1    g629(.A(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n567_), .B2(KEYINPUT60), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n808_), .B(new_n832_), .C1(KEYINPUT60), .C2(new_n831_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n822_), .A2(new_n826_), .A3(new_n567_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n831_), .ZN(G1341gat));
  NAND3_X1  g634(.A1(new_n808_), .A2(new_n226_), .A3(new_n581_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n822_), .A2(new_n826_), .A3(new_n635_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n226_), .ZN(G1342gat));
  INV_X1    g637(.A(new_n605_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n808_), .A2(new_n224_), .A3(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n822_), .A2(new_n826_), .A3(new_n598_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n224_), .ZN(G1343gat));
  INV_X1    g641(.A(new_n806_), .ZN(new_n843_));
  NOR4_X1   g642(.A1(new_n477_), .A2(new_n444_), .A3(new_n482_), .A4(new_n480_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(KEYINPUT124), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  INV_X1    g645(.A(new_n844_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n806_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n644_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(new_n204_), .ZN(G1344gat));
  AOI21_X1  g649(.A(new_n567_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(new_n205_), .ZN(G1345gat));
  AOI21_X1  g651(.A(new_n635_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n853_), .B(new_n855_), .ZN(G1346gat));
  NAND2_X1  g655(.A1(new_n845_), .A2(new_n848_), .ZN(new_n857_));
  INV_X1    g656(.A(G162gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n839_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n598_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n858_), .ZN(G1347gat));
  NOR3_X1   g660(.A1(new_n488_), .A2(new_n391_), .A3(new_n457_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n825_), .A2(new_n444_), .A3(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G169gat), .B1(new_n863_), .B2(new_n644_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n444_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n757_), .B1(new_n818_), .B2(KEYINPUT121), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n824_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n364_), .A3(new_n514_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n865_), .ZN(new_n871_));
  OAI211_X1 g670(.A(G169gat), .B(new_n871_), .C1(new_n863_), .C2(new_n644_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n866_), .A2(new_n870_), .A3(new_n872_), .ZN(G1348gat));
  OAI21_X1  g672(.A(new_n365_), .B1(new_n863_), .B2(new_n567_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n566_), .A2(G176gat), .A3(new_n862_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n806_), .A2(new_n479_), .A3(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n874_), .A2(new_n875_), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G176gat), .B1(new_n869_), .B2(new_n566_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT126), .B1(new_n880_), .B2(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1349gat));
  INV_X1    g681(.A(KEYINPUT127), .ZN(new_n883_));
  INV_X1    g682(.A(new_n346_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n581_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n863_), .B2(new_n885_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n869_), .A2(KEYINPUT127), .A3(new_n884_), .A4(new_n581_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n843_), .A2(new_n444_), .A3(new_n581_), .A4(new_n862_), .ZN(new_n888_));
  INV_X1    g687(.A(G183gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n886_), .A2(new_n887_), .A3(new_n890_), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n863_), .B2(new_n598_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n869_), .A2(new_n347_), .A3(new_n839_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1351gat));
  NOR3_X1   g693(.A1(new_n477_), .A2(new_n484_), .A3(new_n457_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n843_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n644_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n317_), .ZN(G1352gat));
  AOI211_X1 g697(.A(new_n567_), .B(new_n896_), .C1(new_n304_), .C2(new_n302_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n896_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G204gat), .B1(new_n900_), .B2(new_n566_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1353gat));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AND2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n896_), .A2(new_n635_), .A3(new_n903_), .A4(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n900_), .A2(new_n581_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n903_), .ZN(G1354gat));
  OR3_X1    g706(.A1(new_n896_), .A2(G218gat), .A3(new_n605_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G218gat), .B1(new_n896_), .B2(new_n598_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1355gat));
endmodule


