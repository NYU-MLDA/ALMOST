//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT30), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  INV_X1    g004(.A(G15gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G190gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT77), .B(G183gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT25), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  OR3_X1    g013(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n215_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n221_), .B(KEYINPUT23), .ZN(new_n225_));
  INV_X1    g024(.A(new_n210_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(G190gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G169gat), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n214_), .A2(new_n224_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT78), .B1(new_n208_), .B2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(new_n230_), .B2(new_n208_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT31), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n233_), .B(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n223_), .A2(KEYINPUT83), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT83), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n221_), .B(KEYINPUT23), .ZN(new_n241_));
  INV_X1    g040(.A(new_n238_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n229_), .B1(new_n239_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT25), .B(G183gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n209_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n241_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(new_n220_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G211gat), .B(G218gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(KEYINPUT80), .A2(G204gat), .ZN(new_n252_));
  INV_X1    g051(.A(G197gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(KEYINPUT80), .A2(G204gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(G197gat), .B2(G204gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n251_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G197gat), .A2(G204gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n259_), .A2(new_n260_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n250_), .A2(new_n256_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n249_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G226gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n258_), .A2(new_n261_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n230_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n267_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT92), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT92), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n267_), .A2(new_n273_), .A3(new_n276_), .A4(new_n270_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT20), .B1(new_n230_), .B2(new_n272_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n266_), .B1(new_n249_), .B2(KEYINPUT91), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n244_), .B(new_n280_), .C1(new_n220_), .C2(new_n247_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n275_), .B(new_n277_), .C1(new_n282_), .C2(new_n270_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G8gat), .B(G36gat), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n291_), .A3(new_n289_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n283_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n270_), .B1(new_n267_), .B2(new_n273_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT84), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n272_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n270_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n298_), .B1(new_n300_), .B2(new_n278_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n214_), .A2(new_n224_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n227_), .A2(new_n229_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n271_), .B1(new_n304_), .B2(new_n266_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n305_), .A2(KEYINPUT84), .A3(new_n270_), .A4(new_n299_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n297_), .B1(new_n301_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n295_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n296_), .A2(KEYINPUT27), .A3(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n311_));
  NOR2_X1   g110(.A1(new_n307_), .A2(new_n308_), .ZN(new_n312_));
  AOI211_X1 g111(.A(new_n295_), .B(new_n297_), .C1(new_n301_), .C2(new_n306_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G78gat), .B(G106gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318_));
  INV_X1    g117(.A(G141gat), .ZN(new_n319_));
  INV_X1    g118(.A(G148gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n321_), .A2(new_n324_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G141gat), .B(G148gat), .Z(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(KEYINPUT1), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n328_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n329_), .A2(KEYINPUT1), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n332_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n337_), .A2(KEYINPUT29), .ZN(new_n338_));
  OAI211_X1 g137(.A(G228gat), .B(G233gat), .C1(new_n338_), .C2(new_n272_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(KEYINPUT29), .ZN(new_n340_));
  INV_X1    g139(.A(G228gat), .ZN(new_n341_));
  INV_X1    g140(.A(G233gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n266_), .B(new_n340_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n317_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n343_), .A3(new_n317_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n337_), .A2(KEYINPUT29), .ZN(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT79), .B(KEYINPUT28), .Z(new_n349_));
  XNOR2_X1  g148(.A(G22gat), .B(G50gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n348_), .B(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n344_), .B2(KEYINPUT81), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n345_), .A2(KEYINPUT81), .A3(new_n346_), .A4(new_n352_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n315_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G1gat), .B(G29gat), .Z(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT89), .B(KEYINPUT0), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n331_), .A2(new_n336_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n236_), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n234_), .B(new_n235_), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n337_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(KEYINPUT4), .A3(new_n368_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT87), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n365_), .A2(new_n236_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n368_), .A2(KEYINPUT87), .A3(KEYINPUT4), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n371_), .B(new_n372_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n370_), .B1(new_n378_), .B2(KEYINPUT88), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT88), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n372_), .A2(new_n371_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT87), .B1(new_n368_), .B2(KEYINPUT4), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n364_), .B1(new_n379_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n378_), .A2(KEYINPUT88), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n381_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n363_), .A4(new_n370_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n237_), .A2(new_n358_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT94), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT32), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n295_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n283_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT93), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n307_), .B1(new_n393_), .B2(new_n295_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT93), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n283_), .A2(new_n398_), .A3(new_n394_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n396_), .A2(new_n390_), .A3(new_n397_), .A4(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n312_), .A2(new_n313_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n379_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n402_), .A2(KEYINPUT33), .A3(new_n363_), .A4(new_n387_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n384_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n366_), .A2(new_n368_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n405_), .A2(KEYINPUT90), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n371_), .B1(new_n405_), .B2(KEYINPUT90), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n404_), .B(new_n364_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n389_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n401_), .A2(new_n403_), .A3(new_n408_), .A4(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n400_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n392_), .B1(new_n412_), .B2(new_n356_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n356_), .A2(new_n389_), .A3(new_n386_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(KEYINPUT96), .A3(new_n314_), .A4(new_n310_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT96), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n315_), .B2(new_n414_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n356_), .B1(new_n400_), .B2(new_n411_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT94), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n413_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n391_), .B1(new_n422_), .B2(new_n237_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G141gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT76), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G169gat), .B(G197gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT74), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G29gat), .B(G36gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G43gat), .B(G50gat), .Z(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G43gat), .B(G50gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G1gat), .B(G8gat), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439_));
  INV_X1    g238(.A(G1gat), .ZN(new_n440_));
  INV_X1    g239(.A(G8gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT14), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n437_), .A2(new_n442_), .A3(new_n439_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n436_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n435_), .A2(new_n445_), .A3(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G229gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n428_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  AOI211_X1 g251(.A(KEYINPUT74), .B(new_n450_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT75), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n435_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n432_), .A2(new_n434_), .A3(new_n455_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n446_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n454_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n457_), .A2(new_n446_), .A3(KEYINPUT75), .A4(new_n458_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n448_), .A2(new_n450_), .ZN(new_n464_));
  OAI221_X1 g263(.A(new_n427_), .B1(new_n452_), .B2(new_n453_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n427_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n452_), .A2(new_n453_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n464_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G120gat), .B(G148gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT5), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G176gat), .B(G204gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT6), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT9), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(G85gat), .A3(G92gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G85gat), .B(G92gat), .Z(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(KEYINPUT9), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT10), .B(G99gat), .Z(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT64), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT10), .B(G99gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT64), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n491_), .A2(new_n492_), .A3(G106gat), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n482_), .B(new_n487_), .C1(new_n490_), .C2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G57gat), .B(G64gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G71gat), .B(G78gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(KEYINPUT11), .ZN(new_n498_));
  INV_X1    g297(.A(new_n496_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n495_), .A2(KEYINPUT11), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n497_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G99gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(new_n489_), .A3(KEYINPUT65), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT7), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n506_), .A2(new_n503_), .A3(new_n489_), .A4(KEYINPUT65), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n482_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT8), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n486_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n508_), .B2(new_n486_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n494_), .B(new_n502_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT12), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n494_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n502_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n510_), .A2(new_n511_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n508_), .A2(new_n486_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT8), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n508_), .A2(new_n509_), .A3(new_n486_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT66), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n494_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n502_), .A2(KEYINPUT67), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n495_), .A2(KEYINPUT11), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT67), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n497_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n525_), .A2(KEYINPUT12), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(KEYINPUT68), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G85gat), .B(G92gat), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n482_), .B(new_n484_), .C1(new_n483_), .C2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n493_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n492_), .B1(new_n491_), .B2(G106gat), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n518_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n521_), .A2(KEYINPUT66), .A3(new_n522_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n533_), .B1(new_n541_), .B2(new_n530_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n517_), .B1(new_n532_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n516_), .B2(new_n512_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n477_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  AOI211_X1 g347(.A(new_n546_), .B(new_n476_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n472_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n517_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT68), .B1(new_n524_), .B2(new_n531_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n541_), .A2(new_n533_), .A3(new_n530_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n544_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n547_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n476_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n545_), .A2(new_n547_), .A3(new_n477_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(KEYINPUT13), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n550_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT34), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n539_), .A2(new_n540_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n459_), .B1(new_n566_), .B2(new_n494_), .ZN(new_n567_));
  OAI22_X1  g366(.A1(new_n514_), .A2(new_n436_), .B1(KEYINPUT35), .B2(new_n563_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n570_));
  INV_X1    g369(.A(new_n514_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(new_n435_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n572_), .B(new_n564_), .C1(new_n459_), .C2(new_n541_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G134gat), .B(G162gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT70), .Z(new_n579_));
  NAND3_X1  g378(.A1(new_n569_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n569_), .A2(new_n573_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n576_), .B(KEYINPUT36), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n580_), .A2(KEYINPUT71), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT71), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n569_), .A2(new_n573_), .A3(new_n584_), .A4(new_n579_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n561_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n582_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n580_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT73), .B1(new_n586_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n580_), .A2(KEYINPUT71), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT37), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT73), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n589_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT16), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n600_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(KEYINPUT67), .A3(KEYINPUT17), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n515_), .A2(new_n446_), .ZN(new_n605_));
  INV_X1    g404(.A(G231gat), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n342_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n460_), .A2(new_n502_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n605_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n604_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n610_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n605_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n601_), .A2(new_n615_), .A3(new_n602_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n604_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n611_), .B1(new_n614_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n597_), .A2(new_n619_), .ZN(new_n620_));
  NOR4_X1   g419(.A1(new_n423_), .A2(new_n471_), .A3(new_n560_), .A4(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n440_), .A3(new_n390_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n587_), .A2(new_n580_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT97), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n423_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n560_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n470_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n619_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n390_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n622_), .A2(new_n623_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n624_), .A2(new_n635_), .A3(new_n636_), .ZN(G1324gat));
  NAND3_X1  g436(.A1(new_n621_), .A2(new_n441_), .A3(new_n315_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n418_), .B(new_n416_), .C1(new_n420_), .C2(KEYINPUT94), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n420_), .A2(KEYINPUT94), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n237_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n391_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(new_n315_), .A3(new_n626_), .A4(new_n632_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G8gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT98), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n648_), .A3(G8gat), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n646_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n647_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n638_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT40), .B(new_n638_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  INV_X1    g455(.A(new_n237_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n621_), .A2(new_n206_), .A3(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n628_), .A2(new_n657_), .A3(new_n632_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n659_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n659_), .B2(G15gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT99), .Z(G1326gat));
  INV_X1    g462(.A(new_n356_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G22gat), .B1(new_n633_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  INV_X1    g465(.A(G22gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n621_), .A2(new_n667_), .A3(new_n356_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1327gat));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n630_), .A2(new_n619_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  INV_X1    g471(.A(new_n597_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n643_), .B2(new_n673_), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT43), .B(new_n597_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n423_), .B2(new_n597_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n643_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n390_), .A3(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G29gat), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n627_), .A2(new_n631_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n560_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n643_), .A2(new_n470_), .A3(new_n686_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n687_), .A2(G29gat), .A3(new_n634_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n670_), .B1(new_n684_), .B2(new_n689_), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT100), .B(new_n688_), .C1(new_n683_), .C2(G29gat), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1328gat));
  XNOR2_X1  g491(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n678_), .A2(new_n315_), .A3(new_n682_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n315_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n696_), .A2(KEYINPUT101), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(KEYINPUT101), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n643_), .A2(new_n470_), .A3(new_n686_), .A4(new_n700_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT45), .Z(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n693_), .B1(new_n695_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n693_), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n705_), .B(new_n702_), .C1(new_n694_), .C2(G36gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1329gat));
  NAND4_X1  g506(.A1(new_n678_), .A2(new_n682_), .A3(G43gat), .A4(new_n657_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n687_), .A2(new_n237_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(G43gat), .B2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n708_), .B(new_n711_), .C1(G43gat), .C2(new_n709_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1330gat));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n678_), .A2(new_n356_), .A3(new_n682_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G50gat), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n687_), .A2(G50gat), .A3(new_n664_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n716_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT104), .B(new_n719_), .C1(new_n717_), .C2(G50gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1331gat));
  NAND2_X1  g522(.A1(new_n643_), .A2(new_n471_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n724_), .A2(new_n629_), .A3(new_n620_), .ZN(new_n725_));
  INV_X1    g524(.A(G57gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n390_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n465_), .A2(new_n619_), .A3(new_n469_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n629_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n628_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n634_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1332gat));
  NOR2_X1   g531(.A1(new_n699_), .A2(G64gat), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n725_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G64gat), .B1(new_n730_), .B2(new_n699_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT48), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT48), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT105), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n740_), .B(new_n734_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n725_), .A2(new_n743_), .A3(new_n657_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G71gat), .B1(new_n730_), .B2(new_n237_), .ZN(new_n745_));
  XOR2_X1   g544(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n745_), .A2(new_n747_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n744_), .B1(new_n748_), .B2(new_n749_), .ZN(G1334gat));
  OAI21_X1  g549(.A(G78gat), .B1(new_n730_), .B2(new_n664_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT50), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n664_), .A2(G78gat), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT107), .Z(new_n754_));
  NAND2_X1  g553(.A1(new_n725_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n724_), .A2(new_n629_), .A3(new_n685_), .ZN(new_n757_));
  INV_X1    g556(.A(G85gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n390_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n629_), .A2(new_n470_), .A3(new_n619_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(new_n634_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n759_), .B1(new_n764_), .B2(new_n758_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT108), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n763_), .B2(new_n699_), .ZN(new_n767_));
  INV_X1    g566(.A(G92gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n757_), .A2(new_n768_), .A3(new_n315_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1337gat));
  AOI21_X1  g569(.A(new_n503_), .B1(new_n762_), .B2(new_n657_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n685_), .A2(new_n629_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n237_), .A2(new_n491_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n643_), .A2(new_n471_), .A3(new_n772_), .A4(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT109), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT111), .B1(new_n771_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(KEYINPUT110), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n774_), .B(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781_));
  AOI211_X1 g580(.A(new_n237_), .B(new_n761_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n780_), .B(new_n781_), .C1(new_n782_), .C2(new_n503_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n776_), .A2(new_n778_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n778_), .B1(new_n776_), .B2(new_n783_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n757_), .A2(new_n489_), .A3(new_n356_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n489_), .B(new_n788_), .C1(new_n762_), .C2(new_n356_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n788_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n681_), .A2(new_n356_), .A3(new_n760_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G106gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n787_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n787_), .C1(new_n789_), .C2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n555_), .B2(KEYINPUT114), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n476_), .B1(new_n543_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n799_), .B2(new_n555_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n804_), .B(new_n517_), .C1(new_n542_), .C2(new_n532_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n798_), .B1(new_n802_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n554_), .A2(new_n800_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n543_), .A2(new_n803_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(KEYINPUT56), .A4(new_n476_), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n471_), .B(new_n549_), .C1(new_n806_), .C2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n427_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n448_), .A2(new_n451_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n463_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n465_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n626_), .C1(new_n810_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n549_), .B1(new_n806_), .B2(new_n809_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n815_), .B1(new_n818_), .B2(new_n470_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n819_), .B2(new_n627_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n814_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n477_), .B1(new_n554_), .B2(new_n800_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT56), .B1(new_n822_), .B2(new_n808_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n802_), .A2(new_n805_), .A3(new_n798_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n558_), .B(new_n821_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n818_), .A2(KEYINPUT58), .A3(new_n821_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n591_), .A3(new_n596_), .A4(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n816_), .B(new_n820_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT58), .B1(new_n818_), .B2(new_n821_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n597_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT115), .B1(new_n833_), .B2(new_n828_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n631_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n728_), .B(new_n837_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n838_), .A2(new_n550_), .A3(new_n559_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n597_), .A2(new_n836_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n836_), .B1(new_n597_), .B2(new_n839_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n835_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n835_), .A2(KEYINPUT116), .A3(new_n844_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n237_), .A2(new_n358_), .A3(new_n634_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n470_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n829_), .A2(new_n820_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n829_), .A2(new_n820_), .A3(KEYINPUT117), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n816_), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n843_), .B1(new_n859_), .B2(new_n631_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NOR4_X1   g660(.A1(new_n237_), .A2(new_n358_), .A3(KEYINPUT59), .A4(new_n634_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n854_), .A2(new_n470_), .A3(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n853_), .B1(new_n864_), .B2(new_n852_), .ZN(G1340gat));
  NOR2_X1   g664(.A1(new_n629_), .A2(KEYINPUT60), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT118), .B(G120gat), .ZN(new_n867_));
  MUX2_X1   g666(.A(KEYINPUT60), .B(new_n866_), .S(new_n867_), .Z(new_n868_));
  NAND4_X1  g667(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .A4(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT119), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n854_), .A2(new_n560_), .A3(new_n863_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n867_), .ZN(G1341gat));
  AND2_X1   g671(.A1(new_n854_), .A2(new_n863_), .ZN(new_n873_));
  INV_X1    g672(.A(G127gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n631_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n850_), .B2(new_n631_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(KEYINPUT120), .B(new_n874_), .C1(new_n850_), .C2(new_n631_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n873_), .A2(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(G1342gat));
  AOI21_X1  g679(.A(G134gat), .B1(new_n851_), .B2(new_n627_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n673_), .A2(G134gat), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT121), .Z(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n873_), .B2(new_n883_), .ZN(G1343gat));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n829_), .A2(new_n830_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n673_), .A2(KEYINPUT115), .A3(new_n828_), .A4(new_n827_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n816_), .A4(new_n820_), .ZN(new_n888_));
  AOI211_X1 g687(.A(new_n846_), .B(new_n843_), .C1(new_n888_), .C2(new_n631_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT116), .B1(new_n835_), .B2(new_n844_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n699_), .A2(new_n237_), .A3(new_n356_), .A4(new_n390_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n885_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n889_), .A2(new_n890_), .A3(KEYINPUT122), .A4(new_n892_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n470_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT123), .B(G141gat), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n470_), .B(new_n897_), .C1(new_n894_), .C2(new_n895_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1344gat));
  OAI21_X1  g700(.A(new_n560_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G148gat), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n320_), .B(new_n560_), .C1(new_n894_), .C2(new_n895_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1345gat));
  OAI21_X1  g704(.A(new_n619_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n907_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n619_), .B(new_n909_), .C1(new_n894_), .C2(new_n895_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1346gat));
  INV_X1    g710(.A(G162gat), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n912_), .B(new_n627_), .C1(new_n894_), .C2(new_n895_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n847_), .A2(new_n848_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT122), .B1(new_n914_), .B2(new_n892_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n891_), .A2(new_n885_), .A3(new_n893_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n597_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n913_), .B1(new_n917_), .B2(new_n912_), .ZN(G1347gat));
  NOR3_X1   g717(.A1(new_n699_), .A2(new_n237_), .A3(new_n390_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n356_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n860_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n470_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT62), .B1(new_n924_), .B2(KEYINPUT22), .ZN(new_n925_));
  OAI21_X1  g724(.A(G169gat), .B1(new_n924_), .B2(KEYINPUT62), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n216_), .B2(new_n925_), .ZN(G1348gat));
  AOI21_X1  g727(.A(G176gat), .B1(new_n923_), .B2(new_n560_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n914_), .A2(new_n356_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n920_), .A2(new_n217_), .A3(new_n629_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(G1349gat));
  NOR2_X1   g731(.A1(new_n631_), .A2(new_n245_), .ZN(new_n933_));
  AOI21_X1  g732(.A(KEYINPUT124), .B1(new_n923_), .B2(new_n933_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n923_), .A2(KEYINPUT124), .A3(new_n933_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n930_), .A2(new_n619_), .A3(new_n919_), .ZN(new_n936_));
  AOI211_X1 g735(.A(new_n934_), .B(new_n935_), .C1(new_n936_), .C2(new_n210_), .ZN(G1350gat));
  NAND2_X1  g736(.A1(new_n923_), .A2(new_n673_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(G190gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n923_), .A2(new_n209_), .A3(new_n627_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1351gat));
  NOR3_X1   g740(.A1(new_n699_), .A2(new_n657_), .A3(new_n414_), .ZN(new_n942_));
  AND3_X1   g741(.A1(new_n847_), .A2(new_n848_), .A3(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n470_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(KEYINPUT125), .B(G197gat), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n944_), .B(new_n945_), .ZN(G1352gat));
  AOI21_X1  g745(.A(G204gat), .B1(new_n943_), .B2(new_n560_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n943_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n629_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n252_), .A2(new_n254_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n947_), .B1(new_n949_), .B2(new_n950_), .ZN(G1353gat));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n847_), .A2(new_n619_), .A3(new_n848_), .A4(new_n942_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n955_));
  INV_X1    g754(.A(G211gat), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n955_), .A2(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n952_), .B1(new_n954_), .B2(new_n957_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n953_), .A2(KEYINPUT126), .A3(new_n955_), .A4(new_n956_), .ZN(new_n959_));
  XOR2_X1   g758(.A(KEYINPUT63), .B(G211gat), .Z(new_n960_));
  AOI22_X1  g759(.A1(new_n958_), .A2(new_n959_), .B1(new_n954_), .B2(new_n960_), .ZN(G1354gat));
  AOI21_X1  g760(.A(G218gat), .B1(new_n943_), .B2(new_n627_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n673_), .A2(G218gat), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(KEYINPUT127), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n962_), .B1(new_n943_), .B2(new_n964_), .ZN(G1355gat));
endmodule


