//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT15), .Z(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n212_), .A2(new_n204_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G229gat), .A2(G233gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n212_), .B(new_n204_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n215_), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n213_), .A2(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G113gat), .B(G141gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G197gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n219_), .A2(new_n223_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  INV_X1    g033(.A(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n238_), .A2(KEYINPUT9), .ZN(new_n239_));
  INV_X1    g038(.A(G85gat), .ZN(new_n240_));
  INV_X1    g039(.A(G92gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(KEYINPUT9), .A3(new_n238_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n233_), .A2(new_n237_), .A3(new_n239_), .A4(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n242_), .A2(new_n238_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT7), .ZN(new_n247_));
  INV_X1    g046(.A(G99gat), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n235_), .A4(KEYINPUT64), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n250_));
  OAI22_X1  g049(.A1(new_n250_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n231_), .A2(new_n232_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n246_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT8), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n249_), .A2(new_n251_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT8), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n246_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n245_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G71gat), .B(G78gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n261_));
  INV_X1    g060(.A(G57gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(G64gat), .ZN(new_n263_));
  INV_X1    g062(.A(G64gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(G57gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n261_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(G57gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(G64gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT11), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n260_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n260_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n228_), .B1(new_n259_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT65), .B1(new_n270_), .B2(new_n272_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n260_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT11), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT11), .B1(new_n267_), .B2(new_n268_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n271_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n256_), .A2(new_n257_), .A3(new_n246_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n257_), .B1(new_n256_), .B2(new_n246_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n244_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(KEYINPUT12), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G230gat), .A2(G233gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n259_), .A2(new_n273_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n274_), .A2(new_n286_), .A3(new_n287_), .A4(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n287_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n259_), .A2(new_n273_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n273_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n285_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n290_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G120gat), .B(G148gat), .ZN(new_n296_));
  INV_X1    g095(.A(G204gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT5), .B(G176gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n295_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT13), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n301_), .B(KEYINPUT67), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT13), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n212_), .B(new_n310_), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT71), .ZN(new_n312_));
  INV_X1    g111(.A(new_n282_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G127gat), .B(G155gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT16), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(G183gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G211gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT17), .ZN(new_n318_));
  OAI22_X1  g117(.A1(new_n312_), .A2(new_n313_), .B1(KEYINPUT72), .B2(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n312_), .A2(new_n313_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n318_), .A2(KEYINPUT72), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n317_), .A2(KEYINPUT17), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n311_), .B(new_n292_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n318_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n204_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n259_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT68), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT35), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G232gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT34), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n205_), .A2(new_n285_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n333_), .A2(new_n330_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n329_), .B(new_n334_), .C1(new_n330_), .C2(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G190gat), .B(G218gat), .ZN(new_n340_));
  INV_X1    g139(.A(G134gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT69), .ZN(new_n343_));
  INV_X1    g142(.A(G162gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n345_), .A2(KEYINPUT36), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(KEYINPUT36), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n339_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n337_), .A2(new_n346_), .A3(new_n338_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT37), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n348_), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n354_), .A2(KEYINPUT70), .A3(new_n346_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT70), .B1(new_n354_), .B2(new_n346_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n339_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n350_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT37), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n326_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n309_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n227_), .B1(new_n361_), .B2(KEYINPUT73), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT76), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT77), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G71gat), .B(G99gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G15gat), .B(G43gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT78), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n367_), .B(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT74), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(KEYINPUT24), .A3(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT25), .B(G183gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT26), .B(G190gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n375_), .B(new_n378_), .C1(KEYINPUT24), .C2(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT23), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT75), .ZN(new_n383_));
  OAI22_X1  g182(.A1(new_n381_), .A2(KEYINPUT75), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G169gat), .ZN(new_n386_));
  INV_X1    g185(.A(G176gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n388_), .A2(new_n372_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n381_), .B1(G183gat), .B2(G190gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT30), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n370_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n393_), .A2(new_n394_), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n395_), .B(new_n396_), .Z(new_n397_));
  XNOR2_X1  g196(.A(G127gat), .B(G134gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G113gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G120gat), .ZN(new_n402_));
  INV_X1    g201(.A(G113gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n400_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G120gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT31), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n397_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n297_), .A2(G197gat), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n410_), .A2(KEYINPUT86), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(KEYINPUT86), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n222_), .A2(G204gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT21), .ZN(new_n415_));
  XOR2_X1   g214(.A(G211gat), .B(G218gat), .Z(new_n416_));
  INV_X1    g215(.A(KEYINPUT21), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n410_), .A2(new_n413_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n417_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n415_), .A2(new_n419_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT87), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G228gat), .A2(G233gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT84), .ZN(new_n428_));
  NAND3_X1  g227(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT83), .Z(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G141gat), .A2(G148gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT82), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n433_), .B2(KEYINPUT3), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(KEYINPUT3), .B2(new_n433_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n428_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n424_), .A2(KEYINPUT1), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n424_), .B1(new_n426_), .B2(KEYINPUT1), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n439_), .B2(new_n438_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G141gat), .B(G148gat), .Z(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT29), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n422_), .A2(new_n423_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n421_), .B1(new_n444_), .B2(KEYINPUT29), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n423_), .B2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n444_), .A2(KEYINPUT29), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G22gat), .B(G50gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n448_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G78gat), .B(G106gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n455_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n409_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G57gat), .B(G85gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G29gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n463_), .B(new_n464_), .Z(new_n465_));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n407_), .A2(new_n466_), .A3(new_n444_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n444_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n407_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n467_), .B1(new_n470_), .B2(new_n466_), .ZN(new_n471_));
  AND2_X1   g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n469_), .A2(new_n472_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n465_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT33), .B(new_n465_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n465_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n470_), .A2(KEYINPUT98), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT98), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n472_), .B1(new_n469_), .B2(new_n481_), .ZN(new_n482_));
  OAI221_X1 g281(.A(new_n479_), .B1(new_n480_), .B2(new_n482_), .C1(new_n472_), .C2(new_n471_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n477_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n371_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n373_), .B1(new_n487_), .B2(KEYINPUT91), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(KEYINPUT91), .B2(new_n487_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n486_), .A2(new_n374_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n381_), .A4(new_n378_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n389_), .B(KEYINPUT93), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G183gat), .A2(G190gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n494_), .B1(new_n495_), .B2(new_n384_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n492_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n421_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n422_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n392_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n500_), .A2(KEYINPUT20), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G226gat), .A2(G233gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT88), .Z(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT19), .Z(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT89), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT94), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G8gat), .B(G36gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT18), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(G64gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(new_n241_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n422_), .A2(new_n392_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n507_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n516_), .A2(KEYINPUT20), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n515_), .B(new_n517_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n510_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n509_), .A2(KEYINPUT94), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n518_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n514_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n519_), .A2(new_n525_), .A3(KEYINPUT95), .ZN(new_n526_));
  OR3_X1    g325(.A1(new_n523_), .A2(KEYINPUT95), .A3(new_n524_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n526_), .A2(KEYINPUT96), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT96), .B1(new_n526_), .B2(new_n527_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n485_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n474_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n479_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT100), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n475_), .A2(KEYINPUT99), .ZN(new_n534_));
  OR3_X1    g333(.A1(new_n531_), .A2(KEYINPUT99), .A3(new_n479_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n496_), .A2(new_n421_), .A3(new_n491_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n515_), .A2(KEYINPUT20), .A3(new_n538_), .ZN(new_n539_));
  OAI22_X1  g338(.A1(new_n504_), .A2(new_n508_), .B1(new_n516_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(KEYINPUT32), .A3(new_n514_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n514_), .A2(KEYINPUT32), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n510_), .A2(new_n542_), .A3(new_n518_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n537_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n460_), .B1(new_n530_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n409_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(new_n458_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n458_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n409_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT27), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n526_), .A2(new_n527_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n540_), .A2(new_n524_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT101), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(KEYINPUT27), .A3(new_n519_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n550_), .A2(new_n556_), .A3(new_n537_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n545_), .A2(new_n557_), .ZN(new_n558_));
  AOI211_X1 g357(.A(new_n362_), .B(new_n558_), .C1(KEYINPUT73), .C2(new_n361_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n207_), .A3(new_n537_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT38), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n558_), .A2(new_n351_), .A3(new_n326_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n308_), .A2(new_n226_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n537_), .ZN(new_n566_));
  OAI21_X1  g365(.A(G1gat), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n559_), .A2(KEYINPUT38), .A3(new_n207_), .A4(new_n537_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n562_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT102), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(G1324gat));
  INV_X1    g370(.A(new_n556_), .ZN(new_n572_));
  OAI21_X1  g371(.A(G8gat), .B1(new_n565_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n559_), .A2(new_n208_), .A3(new_n556_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT40), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n575_), .A2(KEYINPUT40), .A3(new_n576_), .A4(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(G1325gat));
  INV_X1    g382(.A(G15gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n559_), .A2(new_n584_), .A3(new_n409_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n563_), .A2(new_n564_), .A3(new_n409_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT41), .B1(new_n586_), .B2(G15gat), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n585_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT104), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(G1326gat));
  OAI21_X1  g391(.A(G22gat), .B1(new_n565_), .B2(new_n548_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(G22gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n559_), .A2(new_n596_), .A3(new_n458_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(G1327gat));
  INV_X1    g397(.A(new_n351_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n558_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n326_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n308_), .A2(new_n226_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(G29gat), .B1(new_n604_), .B2(new_n537_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n602_), .B(KEYINPUT106), .Z(new_n606_));
  NAND2_X1  g405(.A1(new_n353_), .A2(new_n359_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT43), .B1(new_n558_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT43), .ZN(new_n609_));
  INV_X1    g408(.A(new_n607_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n609_), .B(new_n610_), .C1(new_n545_), .C2(new_n557_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n606_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT44), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n615_), .A2(G29gat), .A3(new_n537_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n606_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n529_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n526_), .A2(new_n527_), .A3(KEYINPUT96), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n484_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n537_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n459_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n572_), .B(new_n566_), .C1(new_n549_), .C2(new_n547_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n609_), .B1(new_n624_), .B2(new_n610_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n611_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT44), .B(new_n617_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT107), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n612_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n605_), .B1(new_n616_), .B2(new_n631_), .ZN(G1328gat));
  INV_X1    g431(.A(KEYINPUT46), .ZN(new_n633_));
  INV_X1    g432(.A(G36gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n556_), .B1(new_n612_), .B2(KEYINPUT44), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n631_), .B2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n603_), .A2(G36gat), .A3(new_n572_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT45), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n633_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT45), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n638_), .B(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n635_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n642_), .B(KEYINPUT46), .C1(new_n643_), .C2(new_n634_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n644_), .ZN(G1329gat));
  INV_X1    g444(.A(KEYINPUT47), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n603_), .A2(new_n546_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n629_), .A2(new_n630_), .ZN(new_n648_));
  OAI211_X1 g447(.A(G43gat), .B(new_n409_), .C1(new_n612_), .C2(KEYINPUT44), .ZN(new_n649_));
  OAI221_X1 g448(.A(new_n646_), .B1(G43gat), .B2(new_n647_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n647_), .A2(G43gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT47), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(G1330gat));
  AOI21_X1  g453(.A(G50gat), .B1(new_n604_), .B2(new_n458_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n615_), .A2(G50gat), .A3(new_n458_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(new_n631_), .ZN(G1331gat));
  NOR2_X1   g456(.A1(new_n309_), .A2(new_n227_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n563_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G57gat), .B1(new_n659_), .B2(new_n566_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n624_), .A2(new_n360_), .A3(new_n658_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n262_), .A3(new_n537_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1332gat));
  NAND2_X1  g462(.A1(new_n556_), .A2(new_n264_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT108), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n563_), .A2(new_n556_), .A3(new_n658_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT48), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(G64gat), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n667_), .B2(G64gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(G1333gat));
  OAI21_X1  g473(.A(G71gat), .B1(new_n659_), .B2(new_n546_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT49), .ZN(new_n676_));
  INV_X1    g475(.A(G71gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n661_), .A2(new_n677_), .A3(new_n409_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1334gat));
  OAI21_X1  g478(.A(G78gat), .B1(new_n659_), .B2(new_n548_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT50), .ZN(new_n681_));
  INV_X1    g480(.A(G78gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n661_), .A2(new_n682_), .A3(new_n458_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1335gat));
  NAND2_X1  g483(.A1(new_n658_), .A2(new_n326_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n600_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n240_), .A3(new_n537_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n608_), .A2(new_n611_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n566_), .A3(new_n685_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n693_), .B2(new_n240_), .ZN(G1336gat));
  NAND3_X1  g493(.A1(new_n689_), .A2(new_n241_), .A3(new_n556_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n692_), .A2(new_n572_), .A3(new_n685_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n241_), .ZN(G1337gat));
  AND2_X1   g496(.A1(new_n234_), .A2(new_n236_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n689_), .A2(new_n698_), .A3(new_n409_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n692_), .A2(new_n546_), .A3(new_n685_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n248_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT51), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT51), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n699_), .B(new_n703_), .C1(new_n248_), .C2(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1338gat));
  NAND3_X1  g504(.A1(new_n689_), .A2(new_n235_), .A3(new_n458_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n691_), .A2(new_n458_), .A3(new_n686_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT52), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G106gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G106gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT53), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n706_), .B(new_n713_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1339gat));
  INV_X1    g514(.A(KEYINPUT57), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n213_), .A2(new_n214_), .A3(new_n218_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n223_), .B1(new_n217_), .B2(new_n215_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n224_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n303_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT55), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n289_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n289_), .B2(new_n723_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT12), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n255_), .A2(new_n258_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(new_n244_), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n729_), .A2(new_n282_), .B1(new_n273_), .B2(new_n259_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n730_), .A2(KEYINPUT55), .A3(new_n287_), .A4(new_n274_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n286_), .A2(new_n288_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n228_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n290_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n731_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n721_), .B1(new_n726_), .B2(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n731_), .A2(new_n735_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n738_), .B(KEYINPUT112), .C1(new_n725_), .C2(new_n724_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n739_), .A4(new_n300_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(new_n300_), .A3(new_n739_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT56), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n740_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n295_), .A2(new_n300_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n227_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n720_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n716_), .B1(new_n750_), .B2(new_n351_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n289_), .A2(new_n723_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT111), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n289_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n736_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n300_), .B1(new_n755_), .B2(KEYINPUT112), .ZN(new_n756_));
  INV_X1    g555(.A(new_n739_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n743_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT113), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n748_), .B1(new_n761_), .B2(new_n740_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT57), .B(new_n599_), .C1(new_n762_), .C2(new_n720_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n740_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n719_), .A2(new_n747_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n764_), .A2(new_n766_), .B1(KEYINPUT114), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(KEYINPUT114), .ZN(new_n769_));
  AOI211_X1 g568(.A(new_n765_), .B(new_n769_), .C1(new_n758_), .C2(new_n740_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n610_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n751_), .A2(new_n763_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n326_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n309_), .A2(new_n360_), .A3(new_n226_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n774_), .B(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n547_), .A2(new_n537_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n572_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n778_), .A2(new_n779_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n226_), .A2(new_n403_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n771_), .A2(KEYINPUT115), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n610_), .B(new_n788_), .C1(new_n768_), .C2(new_n770_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n751_), .A2(new_n763_), .A3(new_n787_), .A4(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n326_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT116), .B1(new_n791_), .B2(new_n777_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n793_), .B(new_n776_), .C1(new_n790_), .C2(new_n326_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n792_), .A2(new_n794_), .A3(new_n781_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT118), .B1(new_n795_), .B2(new_n779_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n777_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n793_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n791_), .A2(KEYINPUT116), .A3(new_n777_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n782_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(KEYINPUT59), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n784_), .B(new_n786_), .C1(new_n796_), .C2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n792_), .A2(new_n794_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT117), .B1(new_n804_), .B2(new_n782_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  NOR4_X1   g605(.A1(new_n792_), .A2(new_n794_), .A3(new_n806_), .A4(new_n781_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n227_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT119), .B1(new_n803_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n795_), .A2(KEYINPUT117), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n800_), .A2(new_n806_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n403_), .B1(new_n813_), .B2(new_n226_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n795_), .A2(KEYINPUT118), .A3(new_n779_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n801_), .B1(new_n800_), .B2(KEYINPUT59), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n783_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n814_), .B(new_n815_), .C1(new_n818_), .C2(new_n786_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n810_), .A2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(KEYINPUT60), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n309_), .B2(G120gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n811_), .A2(new_n812_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n308_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G120gat), .B1(new_n824_), .B2(new_n818_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(KEYINPUT60), .B2(new_n823_), .ZN(G1341gat));
  OAI21_X1  g625(.A(G127gat), .B1(new_n818_), .B2(new_n326_), .ZN(new_n827_));
  OR3_X1    g626(.A1(new_n813_), .A2(G127gat), .A3(new_n326_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1342gat));
  OAI21_X1  g628(.A(G134gat), .B1(new_n818_), .B2(new_n607_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n808_), .A2(new_n341_), .A3(new_n351_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1343gat));
  NAND3_X1  g631(.A1(new_n572_), .A2(new_n537_), .A3(new_n549_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT120), .Z(new_n834_));
  AND2_X1   g633(.A1(new_n804_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n227_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n308_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g638(.A(KEYINPUT61), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n798_), .A2(new_n601_), .A3(new_n834_), .A4(new_n799_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT121), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n804_), .A2(new_n843_), .A3(new_n601_), .A4(new_n834_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n840_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n844_), .A3(new_n840_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G155gat), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n847_), .ZN(new_n849_));
  INV_X1    g648(.A(G155gat), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n849_), .A2(new_n845_), .A3(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n848_), .A2(new_n851_), .ZN(G1346gat));
  AOI21_X1  g651(.A(G162gat), .B1(new_n835_), .B2(new_n351_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n610_), .A2(G162gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT122), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n835_), .B2(new_n855_), .ZN(G1347gat));
  NOR3_X1   g655(.A1(new_n572_), .A2(new_n537_), .A3(new_n546_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n227_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT123), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(new_n548_), .A3(new_n778_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G169gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT62), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n857_), .A2(new_n548_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n778_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n227_), .A2(new_n386_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n862_), .B1(new_n864_), .B2(new_n865_), .ZN(G1348gat));
  NOR3_X1   g665(.A1(new_n792_), .A2(new_n794_), .A3(new_n458_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n867_), .A2(G176gat), .A3(new_n308_), .A4(new_n857_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n387_), .B1(new_n864_), .B2(new_n309_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT124), .ZN(G1349gat));
  NOR3_X1   g670(.A1(new_n864_), .A2(new_n376_), .A3(new_n326_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n867_), .A2(new_n601_), .A3(new_n857_), .ZN(new_n873_));
  INV_X1    g672(.A(G183gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1350gat));
  OAI21_X1  g674(.A(G190gat), .B1(new_n864_), .B2(new_n607_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n351_), .A2(new_n377_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT125), .Z(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(new_n864_), .B2(new_n878_), .ZN(G1351gat));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n880_));
  AND4_X1   g679(.A1(new_n566_), .A2(new_n804_), .A3(new_n556_), .A4(new_n549_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n227_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n882_), .B2(new_n222_), .ZN(new_n883_));
  AOI211_X1 g682(.A(KEYINPUT126), .B(G197gat), .C1(new_n881_), .C2(new_n227_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n222_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(G1352gat));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n308_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g687(.A1(new_n881_), .A2(new_n601_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  AND2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n889_), .B2(new_n890_), .ZN(G1354gat));
  NAND2_X1  g692(.A1(new_n881_), .A2(new_n351_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT127), .B(G218gat), .Z(new_n895_));
  NOR2_X1   g694(.A1(new_n607_), .A2(new_n895_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n894_), .A2(new_n895_), .B1(new_n881_), .B2(new_n896_), .ZN(G1355gat));
endmodule


