//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT85), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT2), .ZN(new_n205_));
  OR3_X1    g004(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n206_), .B(new_n207_), .C1(new_n208_), .C2(new_n203_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n202_), .B1(new_n205_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT86), .ZN(new_n211_));
  INV_X1    g010(.A(new_n204_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(KEYINPUT1), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(KEYINPUT1), .B2(new_n213_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n212_), .B(new_n216_), .C1(G141gat), .C2(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n211_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT87), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT87), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n211_), .A2(new_n220_), .A3(new_n217_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT89), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n221_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT29), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G197gat), .B(G204gat), .Z(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT21), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(KEYINPUT21), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G211gat), .B(G218gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n231_), .A2(new_n232_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(G228gat), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT91), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n228_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n235_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n218_), .A2(KEYINPUT29), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT92), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n218_), .A2(KEYINPUT92), .A3(KEYINPUT29), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n239_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G78gat), .B(G106gat), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n243_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n241_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n251_), .B1(new_n254_), .B2(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G22gat), .B(G50gat), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n225_), .A2(new_n259_), .A3(new_n226_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT88), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT88), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n260_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n258_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n266_), .A3(new_n258_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n256_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n263_), .A2(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n257_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n272_), .A2(new_n268_), .A3(new_n255_), .A4(new_n253_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT101), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G225gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT97), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G127gat), .B(G134gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G113gat), .B(G120gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n222_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n211_), .A2(new_n281_), .A3(new_n217_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT96), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n219_), .A2(new_n282_), .A3(new_n221_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n277_), .B(new_n283_), .C1(new_n287_), .C2(new_n278_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G1gat), .B(G29gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G57gat), .B(G85gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n277_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n285_), .A2(new_n295_), .A3(new_n286_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n288_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n294_), .B1(new_n288_), .B2(new_n296_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n275_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT101), .A3(new_n297_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT27), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT20), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT22), .B(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT93), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT23), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n310_), .A2(new_n311_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n311_), .B2(new_n310_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT81), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n312_), .B2(KEYINPUT23), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT25), .B(G183gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G190gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G169gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n309_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(KEYINPUT24), .A3(new_n306_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n326_), .A2(KEYINPUT24), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n317_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n305_), .B1(new_n331_), .B2(new_n235_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n313_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n334_));
  AOI21_X1  g133(.A(G176gat), .B1(new_n334_), .B2(KEYINPUT22), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G169gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n320_), .B2(new_n314_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n333_), .A2(new_n337_), .A3(KEYINPUT82), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n332_), .B1(new_n342_), .B2(new_n235_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n341_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT82), .B1(new_n333_), .B2(new_n337_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(new_n244_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT20), .B1(new_n331_), .B2(new_n235_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n351_), .A2(new_n345_), .A3(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G8gat), .B(G36gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n347_), .A2(new_n353_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n351_), .A2(new_n345_), .A3(new_n352_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(new_n346_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n304_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n360_), .A3(new_n346_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n351_), .A2(new_n352_), .ZN(new_n365_));
  MUX2_X1   g164(.A(new_n343_), .B(new_n365_), .S(new_n345_), .Z(new_n366_));
  OAI211_X1 g165(.A(KEYINPUT27), .B(new_n364_), .C1(new_n366_), .C2(new_n360_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n274_), .A2(new_n303_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n361_), .A2(new_n371_), .A3(new_n346_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n366_), .B2(new_n371_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n373_), .B1(new_n301_), .B2(new_n297_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT33), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n297_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT95), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n358_), .B1(new_n347_), .B2(new_n353_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n364_), .A2(new_n379_), .A3(KEYINPUT95), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n288_), .A2(new_n296_), .A3(KEYINPUT33), .A4(new_n294_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n376_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n293_), .B1(new_n287_), .B2(new_n295_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT99), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT99), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n386_), .B(new_n293_), .C1(new_n287_), .C2(new_n295_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n295_), .B(new_n283_), .C1(new_n287_), .C2(new_n278_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT100), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n385_), .A2(KEYINPUT100), .A3(new_n387_), .A4(new_n388_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n374_), .B1(new_n383_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n370_), .B1(new_n394_), .B2(new_n274_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G71gat), .B(G99gat), .ZN(new_n396_));
  INV_X1    g195(.A(G43gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n342_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400_));
  INV_X1    g199(.A(G15gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT30), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n342_), .A2(new_n398_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n399_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n399_), .B2(new_n404_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n281_), .B(KEYINPUT31), .Z(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n409_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n414_));
  OR3_X1    g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n395_), .A2(KEYINPUT102), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT102), .B1(new_n395_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n274_), .A2(new_n368_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(new_n417_), .A3(new_n303_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n419_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G29gat), .B(G36gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT71), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G43gat), .B(G50gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n425_), .A2(KEYINPUT71), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(KEYINPUT71), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n427_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G8gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT73), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G15gat), .B(G22gat), .ZN(new_n436_));
  INV_X1    g235(.A(G1gat), .ZN(new_n437_));
  INV_X1    g236(.A(G8gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT14), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n434_), .A2(KEYINPUT73), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n434_), .A2(KEYINPUT73), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n442_), .A2(new_n439_), .A3(new_n436_), .A4(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n433_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G229gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT15), .ZN(new_n450_));
  INV_X1    g249(.A(new_n432_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n427_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n429_), .A2(KEYINPUT15), .A3(new_n432_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n455_), .A2(KEYINPUT77), .A3(new_n445_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT77), .B1(new_n455_), .B2(new_n445_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n449_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n432_), .A2(new_n429_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n448_), .B1(new_n446_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(KEYINPUT76), .B(new_n448_), .C1(new_n446_), .C2(new_n459_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G113gat), .B(G141gat), .Z(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT78), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G169gat), .B(G197gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n458_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n471_), .B(KEYINPUT79), .Z(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n424_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT12), .ZN(new_n475_));
  INV_X1    g274(.A(G85gat), .ZN(new_n476_));
  INV_X1    g275(.A(G92gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT7), .ZN(new_n487_));
  INV_X1    g286(.A(G99gat), .ZN(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n481_), .B1(new_n486_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT8), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n483_), .A2(new_n485_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(new_n491_), .A3(new_n490_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n481_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n479_), .B1(KEYINPUT65), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT65), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n501_), .A2(new_n503_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n504_));
  OR2_X1    g303(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n489_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT64), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n478_), .A2(new_n502_), .A3(KEYINPUT9), .A4(new_n479_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n505_), .A2(KEYINPUT64), .A3(new_n489_), .A4(new_n506_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n504_), .A2(new_n509_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n475_), .B1(new_n499_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT69), .ZN(new_n514_));
  INV_X1    g313(.A(G57gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(G64gat), .ZN(new_n516_));
  INV_X1    g315(.A(G64gat), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(G57gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT11), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n519_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G71gat), .B(G78gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n522_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n517_), .A2(G57gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n515_), .A2(G64gat), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT11), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n529_), .A2(KEYINPUT66), .A3(new_n524_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n521_), .B1(new_n526_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n523_), .A2(new_n525_), .A3(new_n522_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT66), .B1(new_n529_), .B2(new_n524_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n520_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n531_), .A2(KEYINPUT68), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT68), .B1(new_n531_), .B2(new_n534_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n513_), .B(new_n514_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n490_), .A2(new_n491_), .ZN(new_n538_));
  AOI211_X1 g337(.A(KEYINPUT8), .B(new_n480_), .C1(new_n538_), .C2(new_n495_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n497_), .B1(new_n496_), .B2(new_n481_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n512_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT12), .ZN(new_n542_));
  INV_X1    g341(.A(new_n536_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n531_), .A2(KEYINPUT68), .A3(new_n534_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n499_), .A2(new_n512_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT69), .B1(new_n546_), .B2(KEYINPUT12), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n537_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n531_), .A2(new_n534_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(new_n541_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n550_), .B2(new_n546_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT67), .B(new_n552_), .C1(new_n550_), .C2(new_n546_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n554_), .A2(new_n559_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT70), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n548_), .A2(new_n553_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(KEYINPUT70), .A3(new_n564_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n568_), .A2(new_n564_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT13), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT13), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n455_), .A2(new_n541_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT72), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT34), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT35), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OAI22_X1  g385(.A1(new_n541_), .A2(new_n433_), .B1(KEYINPUT35), .B2(new_n582_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n580_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n586_), .B1(new_n580_), .B2(new_n588_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n589_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n594_), .B(new_n596_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT37), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT37), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n445_), .B(new_n603_), .Z(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(new_n549_), .Z(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  OR3_X1    g411(.A1(new_n605_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT74), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n604_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n604_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n602_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n577_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT75), .Z(new_n621_));
  NAND2_X1  g420(.A1(new_n474_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT103), .ZN(new_n623_));
  INV_X1    g422(.A(new_n303_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n437_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT38), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n576_), .A2(new_n471_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n618_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n598_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n424_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n437_), .B1(new_n632_), .B2(new_n624_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n627_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n634_), .B1(new_n626_), .B2(new_n625_), .ZN(G1324gat));
  XNOR2_X1  g434(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n636_));
  INV_X1    g435(.A(new_n632_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G8gat), .B1(new_n637_), .B2(new_n369_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(KEYINPUT39), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(KEYINPUT39), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n623_), .A2(new_n438_), .A3(new_n368_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n636_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n642_), .B(new_n636_), .C1(new_n640_), .C2(new_n639_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n643_), .A2(new_n645_), .ZN(G1325gat));
  NAND3_X1  g445(.A1(new_n623_), .A2(new_n401_), .A3(new_n417_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n401_), .B1(new_n632_), .B2(new_n417_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT41), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1326gat));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n632_), .B2(new_n274_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT42), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n623_), .A2(new_n651_), .A3(new_n274_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1327gat));
  NOR2_X1   g454(.A1(new_n630_), .A2(new_n598_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n474_), .A2(new_n577_), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G29gat), .B1(new_n657_), .B2(new_n624_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n629_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n602_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT43), .B1(new_n424_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n383_), .A2(new_n393_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n374_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n274_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n368_), .B1(new_n270_), .B2(new_n273_), .ZN(new_n669_));
  AOI22_X1  g468(.A1(new_n667_), .A2(new_n668_), .B1(new_n303_), .B2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n664_), .B1(new_n670_), .B2(new_n417_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n395_), .A2(KEYINPUT102), .A3(new_n418_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n422_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n602_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n630_), .B1(new_n663_), .B2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n659_), .B(new_n661_), .C1(new_n676_), .C2(KEYINPUT105), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n673_), .A2(new_n674_), .A3(new_n602_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n673_), .B2(new_n602_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n618_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n660_), .B(KEYINPUT44), .C1(new_n680_), .C2(new_n629_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n677_), .A2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n624_), .A2(G29gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n658_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  INV_X1    g483(.A(G36gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n657_), .A2(new_n685_), .A3(new_n368_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT45), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n369_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n685_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n687_), .B(new_n690_), .C1(new_n688_), .C2(new_n685_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1329gat));
  NAND3_X1  g493(.A1(new_n657_), .A2(new_n397_), .A3(new_n417_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n418_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n397_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT47), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT47), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n699_), .B(new_n695_), .C1(new_n696_), .C2(new_n397_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1330gat));
  AOI21_X1  g500(.A(G50gat), .B1(new_n657_), .B2(new_n274_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n274_), .A2(G50gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n682_), .B2(new_n703_), .ZN(G1331gat));
  NOR4_X1   g503(.A1(new_n424_), .A2(new_n472_), .A3(new_n577_), .A4(new_n631_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(G57gat), .A3(new_n624_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT107), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT107), .ZN(new_n708_));
  INV_X1    g507(.A(new_n471_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n577_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n673_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n619_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n624_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n707_), .A2(new_n708_), .A3(new_n714_), .ZN(G1332gat));
  AOI21_X1  g514(.A(new_n517_), .B1(new_n705_), .B2(new_n368_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n713_), .A2(new_n517_), .A3(new_n368_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT108), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n717_), .A2(new_n721_), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1333gat));
  INV_X1    g522(.A(G71gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n705_), .B2(new_n417_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n713_), .A2(new_n724_), .A3(new_n417_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1334gat));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n705_), .B2(new_n274_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT50), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n713_), .A2(new_n730_), .A3(new_n274_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1335gat));
  NAND2_X1  g533(.A1(new_n676_), .A2(new_n710_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT110), .Z(new_n736_));
  OAI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n303_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n711_), .A2(new_n656_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n476_), .A3(new_n624_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n736_), .B2(new_n369_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n477_), .A3(new_n368_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n735_), .B2(new_n418_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n738_), .A2(new_n417_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n744_), .A2(new_n745_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n746_), .A2(new_n747_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n738_), .A2(new_n489_), .A3(new_n274_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n676_), .A2(new_n274_), .A3(new_n710_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n753_), .B1(new_n752_), .B2(G106gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n751_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  INV_X1    g558(.A(new_n598_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n553_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n549_), .A2(new_n541_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n514_), .B1(new_n762_), .B2(new_n475_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n513_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n761_), .B1(new_n765_), .B2(new_n537_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n550_), .B1(new_n765_), .B2(new_n537_), .ZN(new_n767_));
  OAI22_X1  g566(.A1(KEYINPUT55), .A2(new_n766_), .B1(new_n767_), .B2(new_n551_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n554_), .A2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n563_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(KEYINPUT56), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n471_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n554_), .A2(new_n769_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n766_), .A2(KEYINPUT55), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n775_), .B(new_n776_), .C1(new_n551_), .C2(new_n767_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT112), .B1(new_n777_), .B2(new_n563_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n773_), .B(new_n774_), .C1(new_n778_), .C2(KEYINPUT56), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n458_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n446_), .A2(new_n447_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n468_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n446_), .A2(new_n459_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n782_), .B(new_n783_), .C1(new_n784_), .C2(new_n448_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n572_), .A2(new_n780_), .A3(new_n785_), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n759_), .B(new_n760_), .C1(new_n779_), .C2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n773_), .A2(new_n774_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n772_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n786_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT57), .B1(new_n790_), .B2(new_n598_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n771_), .A2(KEYINPUT56), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n777_), .A2(new_n793_), .A3(new_n563_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n785_), .A2(new_n780_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT58), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(new_n602_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n797_), .A2(new_n798_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n791_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n787_), .B1(new_n804_), .B2(KEYINPUT118), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(KEYINPUT118), .B2(new_n804_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n618_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n577_), .A2(new_n473_), .A3(new_n619_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT54), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n421_), .A2(new_n417_), .A3(new_n624_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n787_), .A2(new_n791_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n800_), .A2(new_n602_), .A3(new_n803_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n800_), .A2(KEYINPUT114), .A3(new_n602_), .A4(new_n803_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n817_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT115), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n817_), .A2(new_n820_), .A3(new_n824_), .A4(new_n821_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n618_), .A3(new_n825_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n826_), .A2(KEYINPUT116), .A3(new_n809_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT116), .B1(new_n826_), .B2(new_n809_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n811_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n816_), .B1(new_n829_), .B2(new_n813_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n826_), .A2(new_n809_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n826_), .A2(KEYINPUT116), .A3(new_n809_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n812_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n815_), .B1(new_n830_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n473_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n471_), .A2(G113gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n835_), .B2(new_n840_), .ZN(G1340gat));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842_));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n837_), .B2(new_n576_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(KEYINPUT60), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n846_));
  AOI21_X1  g645(.A(G120gat), .B1(new_n576_), .B2(new_n846_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n835_), .A2(new_n845_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n842_), .B1(new_n844_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n815_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n836_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT117), .B1(new_n835_), .B2(KEYINPUT59), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n576_), .B(new_n850_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G120gat), .ZN(new_n854_));
  INV_X1    g653(.A(new_n848_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(KEYINPUT119), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n849_), .A2(new_n856_), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n838_), .B2(new_n618_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n618_), .A2(G127gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n835_), .B2(new_n859_), .ZN(G1342gat));
  OAI21_X1  g659(.A(G134gat), .B1(new_n838_), .B2(new_n662_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n598_), .A2(G134gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n835_), .B2(new_n862_), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n827_), .A2(new_n828_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n668_), .A2(new_n417_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n624_), .A3(new_n369_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n864_), .A2(new_n865_), .A3(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n833_), .A2(new_n834_), .A3(new_n868_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT120), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n709_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  XNOR2_X1  g673(.A(KEYINPUT121), .B(G148gat), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n872_), .B2(new_n576_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI211_X1 g677(.A(KEYINPUT122), .B(new_n577_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n875_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n875_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n877_), .A2(new_n879_), .A3(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1345gat));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n872_), .B2(new_n630_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  AOI211_X1 g687(.A(KEYINPUT123), .B(new_n618_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n885_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n885_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n887_), .A2(new_n889_), .A3(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1346gat));
  INV_X1    g693(.A(new_n872_), .ZN(new_n895_));
  OR3_X1    g694(.A1(new_n895_), .A2(G162gat), .A3(new_n598_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G162gat), .B1(new_n895_), .B2(new_n662_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n624_), .A2(new_n369_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n417_), .A3(new_n668_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n810_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n325_), .B1(new_n901_), .B2(new_n709_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(KEYINPUT124), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n901_), .A2(new_n308_), .A3(new_n709_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n902_), .A2(KEYINPUT124), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT62), .B1(new_n902_), .B2(KEYINPUT124), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n905_), .B(new_n906_), .C1(new_n907_), .C2(new_n908_), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n901_), .B2(new_n576_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n827_), .A2(new_n828_), .A3(new_n274_), .ZN(new_n911_));
  AND4_X1   g710(.A1(G176gat), .A2(new_n899_), .A3(new_n417_), .A4(new_n576_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1349gat));
  NAND4_X1  g712(.A1(new_n911_), .A2(new_n417_), .A3(new_n630_), .A4(new_n899_), .ZN(new_n914_));
  INV_X1    g713(.A(G183gat), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n618_), .A2(new_n322_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n914_), .A2(new_n915_), .B1(new_n901_), .B2(new_n917_), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n901_), .A2(new_n323_), .A3(new_n760_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n810_), .A2(new_n662_), .A3(new_n900_), .ZN(new_n920_));
  INV_X1    g719(.A(G190gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(G1351gat));
  AND2_X1   g721(.A1(new_n866_), .A2(new_n899_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n864_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(KEYINPUT125), .B1(new_n864_), .B2(new_n923_), .ZN(new_n927_));
  OAI211_X1 g726(.A(G197gat), .B(new_n709_), .C1(new_n926_), .C2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n929_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n924_), .B(new_n925_), .ZN(new_n932_));
  AOI21_X1  g731(.A(G197gat), .B1(new_n932_), .B2(new_n709_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n930_), .A2(new_n931_), .A3(new_n933_), .ZN(G1352gat));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n576_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g735(.A(KEYINPUT63), .B(G211gat), .C1(new_n932_), .C2(new_n630_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT63), .B(G211gat), .Z(new_n938_));
  AND3_X1   g737(.A1(new_n932_), .A2(new_n630_), .A3(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1354gat));
  AOI21_X1  g739(.A(G218gat), .B1(new_n932_), .B2(new_n760_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n602_), .A2(G218gat), .ZN(new_n942_));
  XOR2_X1   g741(.A(new_n942_), .B(KEYINPUT127), .Z(new_n943_));
  AOI21_X1  g742(.A(new_n941_), .B1(new_n932_), .B2(new_n943_), .ZN(G1355gat));
endmodule


