//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n956_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_, new_n973_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  XOR2_X1   g001(.A(G57gat), .B(G64gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(KEYINPUT70), .A2(G71gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT70), .A2(G71gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G78gat), .ZN(new_n209_));
  INV_X1    g008(.A(G78gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n210_), .A3(new_n207_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n205_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT71), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n203_), .A2(new_n204_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n205_), .A2(new_n215_), .A3(new_n209_), .A4(new_n211_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n213_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(new_n213_), .B2(new_n216_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n202_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(new_n216_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n214_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT72), .A3(new_n217_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n230_));
  INV_X1    g029(.A(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n233_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n234_), .A2(KEYINPUT66), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT66), .B1(new_n234_), .B2(new_n235_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n229_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G85gat), .B(G92gat), .Z(new_n239_));
  OR2_X1    g038(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n228_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n226_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT68), .B1(new_n227_), .B2(new_n228_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n234_), .A2(new_n235_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT69), .A3(new_n239_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT8), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT69), .B1(new_n248_), .B2(new_n239_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n243_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n236_), .A2(new_n237_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n239_), .A2(KEYINPUT9), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G85gat), .A2(G92gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(KEYINPUT9), .B2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT10), .B(G99gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT64), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n256_), .B1(new_n258_), .B2(new_n232_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n253_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n225_), .A2(KEYINPUT12), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n248_), .A2(new_n239_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT8), .A3(new_n249_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n267_), .A2(new_n243_), .B1(new_n253_), .B2(new_n259_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n223_), .A2(new_n217_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n263_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G230gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n262_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n269_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n261_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n269_), .B1(new_n252_), .B2(new_n260_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n272_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G120gat), .B(G148gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT5), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G176gat), .B(G204gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n284_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n285_), .A2(KEYINPUT13), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT13), .B1(new_n285_), .B2(new_n286_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT76), .B(G1gat), .ZN(new_n290_));
  INV_X1    g089(.A(G8gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT14), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G8gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n294_), .B(KEYINPUT77), .ZN(new_n299_));
  INV_X1    g098(.A(new_n297_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G29gat), .B(G36gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT73), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G43gat), .B(G50gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n298_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n308_));
  OAI211_X1 g107(.A(G229gat), .B(G233gat), .C1(new_n307_), .C2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n298_), .A2(new_n301_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT74), .B(KEYINPUT15), .Z(new_n313_));
  NAND2_X1  g112(.A1(new_n305_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n304_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n303_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n310_), .B(new_n306_), .C1(new_n312_), .C2(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n309_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G113gat), .B(G141gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G169gat), .B(G197gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  OR2_X1    g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n309_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n309_), .A2(new_n320_), .A3(KEYINPUT81), .A4(new_n324_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n289_), .A2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(G231gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n311_), .B(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n334_), .A2(new_n225_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G127gat), .B(G155gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(G183gat), .B(G211gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT17), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n334_), .B2(new_n225_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n335_), .A2(KEYINPUT79), .A3(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n334_), .B(new_n275_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n340_), .A2(KEYINPUT17), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n341_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n332_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G127gat), .B(G134gat), .Z(new_n354_));
  XOR2_X1   g153(.A(G113gat), .B(G120gat), .Z(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G169gat), .ZN(new_n358_));
  INV_X1    g157(.A(G176gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT83), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n362_), .A3(new_n359_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(G183gat), .ZN(new_n365_));
  INV_X1    g164(.A(G190gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT23), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(G183gat), .A3(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT25), .B(G183gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT26), .B(G190gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT24), .A3(new_n374_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n379_), .A2(KEYINPUT24), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n367_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n369_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n368_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  OAI22_X1  g186(.A1(new_n364_), .A2(new_n375_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n389_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(KEYINPUT84), .A3(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G71gat), .B(G99gat), .ZN(new_n394_));
  INV_X1    g193(.A(G43gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(G15gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n396_), .B(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n393_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n403_));
  INV_X1    g202(.A(new_n392_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(new_n390_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n400_), .B1(new_n405_), .B2(new_n393_), .ZN(new_n406_));
  OR3_X1    g205(.A1(new_n402_), .A2(new_n406_), .A3(KEYINPUT31), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT31), .B1(new_n402_), .B2(new_n406_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n357_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(new_n356_), .A3(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n370_), .ZN(new_n418_));
  OR2_X1    g217(.A1(G197gat), .A2(G204gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G197gat), .A2(G204gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT21), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G211gat), .B(G218gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G211gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(G218gat), .ZN(new_n427_));
  INV_X1    g226(.A(G218gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(G211gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT93), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n422_), .A2(new_n425_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n425_), .A2(new_n430_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n419_), .A2(new_n420_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT21), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n432_), .A2(new_n421_), .A3(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n374_), .B(new_n360_), .C1(new_n387_), .C2(new_n371_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n418_), .A2(new_n431_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n431_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n388_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n438_), .A2(new_n440_), .A3(KEYINPUT20), .A4(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT95), .ZN(new_n445_));
  INV_X1    g244(.A(new_n443_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT20), .B1(new_n388_), .B2(new_n439_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n437_), .A2(new_n418_), .B1(new_n431_), .B2(new_n436_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n445_), .B(new_n446_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n360_), .A2(new_n374_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n385_), .A2(new_n386_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n367_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n453_), .B2(new_n372_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n367_), .A2(new_n369_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n382_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n439_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n417_), .A2(new_n453_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n361_), .A2(new_n374_), .A3(new_n373_), .A4(new_n363_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n431_), .A3(new_n459_), .A4(new_n436_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n460_), .A3(KEYINPUT20), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n445_), .B1(new_n461_), .B2(new_n446_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n444_), .B1(new_n450_), .B2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G8gat), .B(G36gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G64gat), .B(G92gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n463_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n468_), .B(new_n444_), .C1(new_n450_), .C2(new_n462_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT97), .A3(new_n471_), .ZN(new_n472_));
  OR3_X1    g271(.A1(new_n463_), .A2(KEYINPUT97), .A3(new_n469_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT27), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT103), .B(KEYINPUT20), .Z(new_n476_));
  NAND3_X1  g275(.A1(new_n438_), .A2(new_n440_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n446_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n446_), .B2(new_n461_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n469_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n471_), .A2(new_n480_), .A3(KEYINPUT27), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(new_n210_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(new_n232_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n488_));
  NOR2_X1   g287(.A1(G155gat), .A2(G162gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT86), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G155gat), .A2(G162gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n494_));
  NOR4_X1   g293(.A1(new_n494_), .A2(KEYINPUT87), .A3(G141gat), .A4(G148gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(G141gat), .A2(G148gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT3), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G141gat), .A2(G148gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT2), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n499_), .A2(KEYINPUT88), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT88), .B1(new_n499_), .B2(new_n500_), .ZN(new_n502_));
  OAI22_X1  g301(.A1(new_n495_), .A2(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n493_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G141gat), .ZN(new_n508_));
  INV_X1    g307(.A(G148gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n497_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n494_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n496_), .A2(new_n497_), .A3(KEYINPUT3), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n499_), .A2(new_n500_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n499_), .A2(KEYINPUT88), .A3(new_n500_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n504_), .B(KEYINPUT89), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n513_), .A2(new_n518_), .A3(new_n519_), .A4(KEYINPUT90), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n492_), .B1(new_n507_), .B2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n491_), .B(KEYINPUT1), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n490_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n496_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n499_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n528_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n488_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n488_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n487_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n439_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G22gat), .B(G50gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n533_), .A2(new_n536_), .A3(new_n487_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n542_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n545_), .B2(new_n537_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n416_), .A2(new_n483_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n492_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n511_), .A2(new_n512_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT90), .B1(new_n550_), .B2(new_n519_), .ZN(new_n551_));
  AND4_X1   g350(.A1(KEYINPUT90), .A2(new_n513_), .A3(new_n518_), .A4(new_n519_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n549_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(new_n357_), .A3(new_n525_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n356_), .B1(new_n521_), .B2(new_n526_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT98), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n525_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT98), .A3(new_n356_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT4), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G225gat), .A2(G233gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n555_), .A2(KEYINPUT4), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT100), .ZN(new_n567_));
  XOR2_X1   g366(.A(G1gat), .B(G29gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT99), .B(G85gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT0), .B(G57gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n563_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n565_), .A2(new_n567_), .A3(new_n573_), .A4(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT104), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n574_), .B(KEYINPUT100), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n580_), .A2(KEYINPUT104), .A3(new_n573_), .A4(new_n565_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n565_), .A2(new_n567_), .A3(new_n576_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n572_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT105), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT105), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n583_), .A2(new_n586_), .A3(new_n572_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n582_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n548_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT106), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n475_), .A2(new_n543_), .A3(new_n546_), .A4(new_n481_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n585_), .A2(new_n587_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n591_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(KEYINPUT106), .A4(new_n582_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n463_), .B1(KEYINPUT32), .B2(new_n468_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n479_), .A2(KEYINPUT32), .A3(new_n468_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n472_), .A2(new_n473_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT102), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n562_), .B1(new_n560_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n600_), .B2(new_n560_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n561_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n572_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n577_), .B2(KEYINPUT101), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n577_), .A2(KEYINPUT101), .A3(new_n606_), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n588_), .A2(new_n598_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n547_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n592_), .B(new_n595_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n416_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n589_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT34), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n252_), .A2(new_n260_), .A3(new_n305_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n319_), .B1(new_n252_), .B2(new_n260_), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT35), .B(new_n616_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n319_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n261_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n268_), .A2(new_n305_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .A4(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n619_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n629_), .A2(KEYINPUT36), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n629_), .B(KEYINPUT36), .Z(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n626_), .B2(KEYINPUT75), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT75), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n619_), .A2(new_n625_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n631_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n614_), .A2(KEYINPUT108), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT108), .B1(new_n614_), .B2(new_n639_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n353_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n588_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n331_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT80), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n347_), .A2(new_n647_), .A3(new_n350_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n637_), .A2(KEYINPUT37), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT37), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n653_), .B(new_n631_), .C1(new_n626_), .C2(new_n632_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(new_n289_), .A3(new_n655_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n614_), .A2(new_n646_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n588_), .A3(new_n290_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT38), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n645_), .A2(new_n659_), .ZN(G1324gat));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n291_), .A3(new_n482_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n642_), .A2(new_n482_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(G8gat), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT39), .B(new_n291_), .C1(new_n642_), .C2(new_n482_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT40), .B(new_n661_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1325gat));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n642_), .A2(new_n416_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(G15gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n672_), .B2(G15gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n671_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n676_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n678_), .A2(KEYINPUT41), .A3(new_n674_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n657_), .A2(new_n398_), .A3(new_n416_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n679_), .A3(new_n680_), .ZN(G1326gat));
  INV_X1    g480(.A(G22gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n657_), .A2(new_n682_), .A3(new_n611_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G22gat), .B1(new_n643_), .B2(new_n547_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT42), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(KEYINPUT42), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(G1327gat));
  NAND2_X1  g486(.A1(new_n595_), .A2(new_n592_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n588_), .A2(new_n598_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n608_), .A2(new_n609_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n611_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n613_), .B1(new_n688_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n589_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n650_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n648_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n639_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n694_), .A2(new_n331_), .A3(new_n289_), .A4(new_n698_), .ZN(new_n699_));
  OR3_X1    g498(.A1(new_n699_), .A2(G29gat), .A3(new_n644_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n655_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(KEYINPUT111), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n704_), .B(KEYINPUT43), .C1(new_n614_), .C2(new_n655_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  OR3_X1    g505(.A1(new_n332_), .A2(KEYINPUT110), .A3(new_n651_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT110), .B1(new_n332_), .B2(new_n651_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n706_), .A2(KEYINPUT44), .A3(new_n710_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n588_), .A3(new_n714_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n715_), .A2(KEYINPUT112), .A3(G29gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT112), .B1(new_n715_), .B2(G29gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n700_), .B1(new_n716_), .B2(new_n717_), .ZN(G1328gat));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  INV_X1    g518(.A(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n706_), .B2(new_n710_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n712_), .B(new_n709_), .C1(new_n703_), .C2(new_n705_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n720_), .B1(new_n723_), .B2(new_n482_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n699_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n720_), .A3(new_n482_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT45), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n719_), .B1(new_n724_), .B2(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n721_), .A2(new_n722_), .A3(new_n483_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT46), .B(new_n727_), .C1(new_n730_), .C2(new_n720_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1329gat));
  NOR4_X1   g531(.A1(new_n721_), .A2(new_n722_), .A3(new_n395_), .A4(new_n613_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n395_), .B1(new_n699_), .B2(new_n613_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT113), .Z(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT47), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n723_), .A2(G43gat), .A3(new_n416_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n735_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(new_n740_), .ZN(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n725_), .B2(new_n611_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n611_), .A2(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n723_), .B2(new_n743_), .ZN(G1331gat));
  OR2_X1    g543(.A1(new_n652_), .A2(new_n654_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(new_n696_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n289_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT114), .Z(new_n749_));
  NAND2_X1  g548(.A1(new_n694_), .A2(new_n646_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G57gat), .B1(new_n753_), .B2(new_n588_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n640_), .A2(new_n641_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n755_), .A2(new_n646_), .A3(new_n747_), .A4(new_n651_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n588_), .B2(KEYINPUT115), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(KEYINPUT115), .B2(new_n758_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n754_), .B1(new_n757_), .B2(new_n760_), .ZN(G1332gat));
  OR3_X1    g560(.A1(new_n752_), .A2(G64gat), .A3(new_n483_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n757_), .A2(new_n482_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(G64gat), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G64gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(G1333gat));
  INV_X1    g566(.A(G71gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n753_), .A2(new_n768_), .A3(new_n416_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n757_), .A2(new_n416_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G71gat), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT49), .B(new_n768_), .C1(new_n757_), .C2(new_n416_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1334gat));
  NAND3_X1  g573(.A1(new_n753_), .A2(new_n210_), .A3(new_n611_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n757_), .A2(new_n611_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(G78gat), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT50), .B(new_n210_), .C1(new_n757_), .C2(new_n611_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1335gat));
  NAND3_X1  g579(.A1(new_n747_), .A2(new_n646_), .A3(new_n696_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n644_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n750_), .A2(new_n289_), .A3(new_n697_), .ZN(new_n785_));
  INV_X1    g584(.A(G85gat), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(new_n588_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(G1336gat));
  OAI21_X1  g587(.A(G92gat), .B1(new_n783_), .B2(new_n483_), .ZN(new_n789_));
  INV_X1    g588(.A(G92gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n785_), .A2(new_n790_), .A3(new_n482_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1337gat));
  AOI21_X1  g591(.A(new_n231_), .B1(new_n782_), .B2(new_n416_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n785_), .A2(new_n416_), .A3(new_n258_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g596(.A1(new_n785_), .A2(new_n232_), .A3(new_n611_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n782_), .A2(new_n611_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(G106gat), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n232_), .B(new_n799_), .C1(new_n782_), .C2(new_n611_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n798_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT53), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n798_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n306_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n310_), .B1(new_n810_), .B2(KEYINPUT118), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(KEYINPUT118), .B2(new_n810_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n307_), .A2(new_n308_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n324_), .B1(new_n813_), .B2(new_n310_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n330_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n220_), .A2(new_n224_), .A3(KEYINPUT12), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n277_), .A2(KEYINPUT12), .B1(new_n818_), .B2(new_n268_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n272_), .B1(new_n819_), .B2(new_n276_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n271_), .B1(new_n261_), .B2(new_n275_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n819_), .B2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n262_), .A2(KEYINPUT55), .A3(new_n270_), .A4(new_n273_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n820_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n283_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n283_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n331_), .A2(new_n286_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n817_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n809_), .B1(new_n833_), .B2(new_n639_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT107), .B(new_n631_), .C1(new_n636_), .C2(new_n634_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n634_), .A2(new_n636_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n631_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n638_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n831_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n840_), .B(KEYINPUT119), .C1(new_n841_), .C2(new_n817_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n834_), .A2(new_n835_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n816_), .B1(new_n279_), .B2(new_n284_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n283_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n845_), .A2(KEYINPUT120), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n829_), .B1(new_n845_), .B2(KEYINPUT120), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT58), .B(new_n844_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n850_), .A2(KEYINPUT121), .A3(new_n745_), .A4(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n840_), .B(KEYINPUT57), .C1(new_n841_), .C2(new_n817_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n843_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(new_n745_), .A3(new_n851_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n351_), .B1(new_n854_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n746_), .A2(new_n859_), .A3(new_n646_), .A4(new_n289_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT54), .B1(new_n656_), .B2(new_n331_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n858_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n858_), .A2(KEYINPUT122), .A3(new_n863_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n548_), .A2(new_n644_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G113gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n331_), .ZN(new_n872_));
  OR3_X1    g671(.A1(new_n548_), .A2(KEYINPUT59), .A3(new_n644_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n843_), .A2(KEYINPUT123), .A3(new_n855_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n853_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT123), .B1(new_n843_), .B2(new_n855_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n696_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n873_), .B1(new_n877_), .B2(new_n863_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n646_), .B(new_n878_), .C1(new_n869_), .C2(KEYINPUT59), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n872_), .B1(new_n879_), .B2(new_n871_), .ZN(G1340gat));
  INV_X1    g679(.A(G120gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n289_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n870_), .B(new_n882_), .C1(KEYINPUT60), .C2(new_n881_), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n289_), .B(new_n878_), .C1(new_n869_), .C2(KEYINPUT59), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n881_), .ZN(G1341gat));
  INV_X1    g684(.A(G127gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n870_), .A2(new_n886_), .A3(new_n651_), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n351_), .B(new_n878_), .C1(new_n869_), .C2(KEYINPUT59), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n886_), .ZN(G1342gat));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n870_), .A2(new_n890_), .A3(new_n639_), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n655_), .B(new_n878_), .C1(new_n869_), .C2(KEYINPUT59), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n890_), .ZN(G1343gat));
  NAND2_X1  g692(.A1(new_n855_), .A2(new_n856_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n894_), .A2(new_n852_), .A3(new_n843_), .A4(new_n853_), .ZN(new_n895_));
  AOI211_X1 g694(.A(new_n865_), .B(new_n862_), .C1(new_n895_), .C2(new_n351_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT122), .B1(new_n858_), .B2(new_n863_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n416_), .A2(new_n547_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n588_), .A3(new_n483_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n331_), .A3(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g702(.A1(new_n898_), .A2(new_n747_), .A3(new_n901_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g704(.A1(new_n898_), .A2(new_n651_), .A3(new_n901_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1346gat));
  INV_X1    g707(.A(G162gat), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n898_), .A2(new_n909_), .A3(new_n639_), .A4(new_n901_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n866_), .A2(new_n867_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n911_), .A2(new_n655_), .A3(new_n900_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n912_), .B2(new_n909_), .ZN(G1347gat));
  NAND2_X1  g712(.A1(new_n877_), .A2(new_n863_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n416_), .A2(new_n547_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n915_), .A2(new_n588_), .A3(new_n483_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n331_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n917_), .A2(new_n918_), .A3(G169gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n917_), .B2(G169gat), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n916_), .ZN(new_n923_));
  AOI211_X1 g722(.A(KEYINPUT124), .B(new_n923_), .C1(new_n877_), .C2(new_n863_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n331_), .A2(new_n358_), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT125), .Z(new_n927_));
  OAI22_X1  g726(.A1(new_n919_), .A2(new_n920_), .B1(new_n925_), .B2(new_n927_), .ZN(G1348gat));
  OAI21_X1  g727(.A(new_n747_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n923_), .A2(new_n359_), .A3(new_n289_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n929_), .A2(new_n359_), .B1(new_n898_), .B2(new_n930_), .ZN(G1349gat));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n351_), .A2(new_n376_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n843_), .A2(new_n855_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n937_), .A2(new_n853_), .A3(new_n874_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n862_), .B1(new_n938_), .B2(new_n696_), .ZN(new_n939_));
  OAI21_X1  g738(.A(KEYINPUT124), .B1(new_n939_), .B2(new_n923_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n914_), .A2(new_n921_), .A3(new_n916_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n934_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n923_), .A2(new_n696_), .ZN(new_n943_));
  AOI21_X1  g742(.A(G183gat), .B1(new_n898_), .B2(new_n943_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n932_), .B1(new_n942_), .B2(new_n944_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n933_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n943_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n365_), .B1(new_n911_), .B2(new_n947_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n946_), .A2(KEYINPUT126), .A3(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n945_), .A2(new_n949_), .ZN(G1350gat));
  AOI21_X1  g749(.A(new_n655_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n639_), .A2(new_n377_), .ZN(new_n952_));
  OAI22_X1  g751(.A1(new_n951_), .A2(new_n366_), .B1(new_n925_), .B2(new_n952_), .ZN(G1351gat));
  NAND3_X1  g752(.A1(new_n899_), .A2(new_n644_), .A3(new_n482_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n898_), .A2(new_n331_), .A3(new_n955_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g756(.A1(new_n911_), .A2(new_n954_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n747_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(G204gat), .ZN(new_n960_));
  INV_X1    g759(.A(G204gat), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n958_), .A2(new_n961_), .A3(new_n747_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n960_), .A2(new_n962_), .ZN(G1353gat));
  INV_X1    g762(.A(new_n351_), .ZN(new_n964_));
  XOR2_X1   g763(.A(KEYINPUT63), .B(G211gat), .Z(new_n965_));
  NAND3_X1  g764(.A1(new_n958_), .A2(new_n964_), .A3(new_n965_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n898_), .A2(new_n964_), .A3(new_n955_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n967_), .A2(new_n968_), .A3(new_n426_), .ZN(new_n969_));
  AND2_X1   g768(.A1(new_n966_), .A2(new_n969_), .ZN(G1354gat));
  NAND2_X1  g769(.A1(new_n958_), .A2(new_n639_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n655_), .A2(new_n428_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(KEYINPUT127), .ZN(new_n973_));
  AOI22_X1  g772(.A1(new_n971_), .A2(new_n428_), .B1(new_n958_), .B2(new_n973_), .ZN(G1355gat));
endmodule


