//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT3), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT2), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT85), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT85), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n208_), .A3(new_n205_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT86), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT87), .ZN(new_n217_));
  OR3_X1    g016(.A1(new_n212_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT84), .B1(new_n212_), .B2(KEYINPUT1), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .A4(new_n211_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n202_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n204_), .A3(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n216_), .A2(new_n217_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n214_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n223_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT87), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G127gat), .B(G134gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT83), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n228_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n225_), .A2(new_n226_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n231_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT97), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n234_), .A2(new_n241_), .A3(KEYINPUT4), .A4(new_n236_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT97), .B1(new_n234_), .B2(KEYINPUT4), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n232_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n236_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n242_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n240_), .B1(new_n248_), .B2(new_n239_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G1gat), .B(G29gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G85gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT0), .B(G57gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G64gat), .B(G92gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(G8gat), .B(G36gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT23), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(G183gat), .A3(G190gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT81), .ZN(new_n265_));
  INV_X1    g064(.A(G183gat), .ZN(new_n266_));
  INV_X1    g065(.A(G190gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT23), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n266_), .A2(KEYINPUT25), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(KEYINPUT25), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n275_));
  INV_X1    g074(.A(G169gat), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G169gat), .B(G176gat), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n275_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n269_), .A2(new_n274_), .A3(new_n279_), .A4(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT93), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n268_), .A2(new_n264_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(G183gat), .B2(G190gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n276_), .A2(new_n277_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT22), .B(G169gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n277_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT94), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n293_), .A2(KEYINPUT89), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n295_), .B1(new_n294_), .B2(new_n293_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n292_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT95), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n301_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n269_), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n289_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n285_), .B1(KEYINPUT24), .B2(new_n278_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(KEYINPUT24), .B2(new_n280_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n271_), .B(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT80), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n311_), .A2(KEYINPUT80), .A3(new_n270_), .A4(new_n273_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n309_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n305_), .A2(new_n307_), .A3(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n317_), .A2(KEYINPUT20), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n292_), .A2(KEYINPUT95), .A3(new_n301_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n304_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT19), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n284_), .A2(new_n305_), .A3(new_n291_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n316_), .A2(new_n307_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n301_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n324_), .A2(KEYINPUT20), .A3(new_n325_), .A4(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n262_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  AOI211_X1 g129(.A(new_n261_), .B(new_n330_), .C1(new_n320_), .C2(new_n322_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n253_), .B1(new_n248_), .B2(new_n238_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(new_n238_), .B2(new_n237_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n249_), .B(new_n253_), .C1(KEYINPUT98), .C2(KEYINPUT33), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n256_), .A2(new_n332_), .A3(new_n334_), .A4(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n253_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n241_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n237_), .B2(new_n246_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n238_), .B1(new_n339_), .B2(new_n242_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n337_), .B1(new_n340_), .B2(new_n240_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n254_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n323_), .A2(new_n328_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n262_), .A2(KEYINPUT32), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n320_), .A2(new_n322_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n282_), .A2(new_n290_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT99), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n305_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(KEYINPUT100), .A3(KEYINPUT20), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n327_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT100), .B1(new_n349_), .B2(KEYINPUT20), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n322_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n346_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n344_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n342_), .A2(new_n345_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n336_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI211_X1 g158(.A(new_n359_), .B(new_n305_), .C1(new_n228_), .C2(KEYINPUT29), .ZN(new_n360_));
  XOR2_X1   g159(.A(G78gat), .B(G106gat), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT29), .B1(new_n225_), .B2(new_n226_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n358_), .B1(new_n363_), .B2(new_n301_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n228_), .B2(KEYINPUT29), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G22gat), .B(G50gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369_));
  INV_X1    g168(.A(new_n366_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n224_), .A2(new_n227_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n368_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n365_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT90), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n362_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n374_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT90), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n372_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n228_), .A2(KEYINPUT29), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(new_n358_), .A3(new_n301_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n364_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n361_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n377_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n381_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT91), .B1(new_n378_), .B2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n381_), .B(new_n362_), .C1(new_n364_), .C2(new_n360_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n376_), .A2(new_n385_), .A3(new_n377_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT91), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .A4(new_n375_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n357_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n331_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n320_), .A2(new_n322_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n352_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(new_n327_), .A3(new_n350_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n322_), .B2(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n395_), .B(KEYINPUT27), .C1(new_n399_), .C2(new_n262_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n342_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n394_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G15gat), .B(G43gat), .Z(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  NAND2_X1  g210(.A1(new_n326_), .A2(KEYINPUT30), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n316_), .A2(new_n307_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT82), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n412_), .A2(new_n417_), .A3(new_n414_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n411_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n411_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n232_), .B(KEYINPUT31), .Z(new_n423_));
  NOR3_X1   g222(.A1(new_n419_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n418_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n421_), .B1(new_n426_), .B2(new_n420_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n422_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n425_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n341_), .A2(new_n254_), .A3(new_n430_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(new_n388_), .A3(new_n392_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n400_), .A2(new_n402_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT101), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n432_), .A2(new_n392_), .A3(new_n388_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT101), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n403_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n406_), .A2(new_n431_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT11), .ZN(new_n440_));
  OR2_X1    g239(.A1(G57gat), .A2(G64gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G57gat), .A2(G64gat), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(G57gat), .A2(G64gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G57gat), .A2(G64gat), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n445_), .A2(new_n446_), .A3(KEYINPUT11), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G71gat), .B(G78gat), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n447_), .A2(KEYINPUT67), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450_));
  XOR2_X1   g249(.A(G71gat), .B(G78gat), .Z(new_n451_));
  NAND3_X1  g250(.A1(new_n441_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n444_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT67), .B1(new_n447_), .B2(new_n448_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n452_), .A3(new_n450_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n443_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G231gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G15gat), .B(G22gat), .ZN(new_n461_));
  INV_X1    g260(.A(G1gat), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G8gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n466_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n469_), .B(KEYINPUT76), .Z(new_n470_));
  XNOR2_X1  g269(.A(new_n460_), .B(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G127gat), .B(G155gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G211gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT16), .B(G183gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n471_), .A2(KEYINPUT17), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(KEYINPUT17), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n471_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481_));
  XOR2_X1   g280(.A(G43gat), .B(G50gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(G29gat), .B(G36gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT15), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT64), .ZN(new_n487_));
  AND3_X1   g286(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(KEYINPUT64), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G85gat), .B(G92gat), .Z(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT9), .ZN(new_n498_));
  XOR2_X1   g297(.A(KEYINPUT10), .B(G99gat), .Z(new_n499_));
  INV_X1    g298(.A(G106gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT9), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(G85gat), .A3(G92gat), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n496_), .A2(new_n498_), .A3(new_n501_), .A4(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT8), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n488_), .A2(new_n489_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n500_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT66), .A3(new_n507_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n505_), .B1(new_n516_), .B2(new_n497_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n507_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n497_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n504_), .B1(new_n517_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n486_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT34), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n527_), .A2(KEYINPUT35), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n525_), .B(new_n528_), .C1(new_n484_), .C2(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(KEYINPUT35), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT36), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT73), .B(KEYINPUT74), .Z(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G134gat), .B(G162gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n532_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n531_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT36), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n481_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n545_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(KEYINPUT37), .A3(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n439_), .A2(new_n480_), .A3(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n469_), .A2(new_n484_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n486_), .A2(new_n469_), .B1(KEYINPUT77), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n469_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n485_), .A2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n552_), .B1(KEYINPUT77), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n469_), .B(new_n484_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n557_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT78), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n557_), .A2(new_n560_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n563_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n567_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT68), .ZN(new_n571_));
  INV_X1    g370(.A(new_n504_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n516_), .A2(new_n497_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT8), .ZN(new_n574_));
  INV_X1    g373(.A(new_n519_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n497_), .A3(new_n521_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n572_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n571_), .B1(new_n577_), .B2(new_n458_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT12), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n458_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n454_), .A2(new_n457_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n524_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n571_), .A3(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .A4(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n583_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n580_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G176gat), .B(G204gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(G120gat), .B(G148gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n586_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT71), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n586_), .A2(new_n589_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(KEYINPUT70), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(KEYINPUT70), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n596_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT13), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n599_), .B(KEYINPUT70), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT13), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n596_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT72), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n550_), .A2(new_n570_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(new_n462_), .A3(new_n342_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n544_), .A2(new_n545_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n439_), .A2(new_n613_), .A3(new_n480_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n607_), .A2(new_n570_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n342_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n609_), .A2(KEYINPUT38), .A3(new_n462_), .A4(new_n342_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n612_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(G1324gat));
  NAND3_X1  g421(.A1(new_n614_), .A2(new_n615_), .A3(new_n434_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(G8gat), .A3(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n623_), .A2(G8gat), .A3(new_n628_), .A4(new_n624_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n550_), .A2(new_n570_), .A3(new_n608_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n434_), .A2(new_n463_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n630_), .A2(KEYINPUT103), .A3(new_n631_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n627_), .B(new_n629_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  OAI21_X1  g437(.A(G15gat), .B1(new_n616_), .B2(new_n431_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT41), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n630_), .A2(G15gat), .A3(new_n431_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1326gat));
  XOR2_X1   g441(.A(new_n393_), .B(KEYINPUT106), .Z(new_n643_));
  OAI21_X1  g442(.A(G22gat), .B1(new_n616_), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT42), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n643_), .A2(G22gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n630_), .B2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(new_n613_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n439_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n615_), .A3(new_n480_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n342_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n546_), .A2(new_n548_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n549_), .B2(KEYINPUT107), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n439_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT107), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT43), .B1(new_n653_), .B2(new_n657_), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n357_), .A2(new_n393_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n437_), .B1(new_n436_), .B2(new_n403_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n433_), .A2(new_n434_), .A3(KEYINPUT101), .ZN(new_n661_));
  OAI22_X1  g460(.A1(new_n659_), .A2(new_n430_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n658_), .B1(new_n662_), .B2(new_n549_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n615_), .B(new_n480_), .C1(new_n656_), .C2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n655_), .B1(new_n439_), .B2(new_n653_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(new_n658_), .A3(new_n549_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n669_), .A2(KEYINPUT44), .A3(new_n615_), .A4(new_n480_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n666_), .A2(new_n342_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n652_), .B1(new_n671_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n434_), .A3(new_n670_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G36gat), .ZN(new_n674_));
  OR4_X1    g473(.A1(KEYINPUT45), .A2(new_n650_), .A3(G36gat), .A4(new_n403_), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n651_), .A2(new_n676_), .A3(new_n434_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT45), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n674_), .A2(new_n679_), .A3(KEYINPUT46), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  NAND4_X1  g483(.A1(new_n666_), .A2(G43gat), .A3(new_n430_), .A4(new_n670_), .ZN(new_n685_));
  INV_X1    g484(.A(G43gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n650_), .B2(new_n431_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g488(.A(new_n643_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G50gat), .B1(new_n651_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n393_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n666_), .A2(new_n692_), .A3(new_n670_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n693_), .B2(G50gat), .ZN(G1331gat));
  NOR2_X1   g493(.A1(new_n608_), .A2(new_n570_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n614_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(G57gat), .A3(new_n342_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT108), .Z(new_n698_));
  NOR2_X1   g497(.A1(new_n607_), .A2(new_n570_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n550_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n342_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n698_), .A2(new_n702_), .ZN(G1332gat));
  INV_X1    g502(.A(G64gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n696_), .B2(new_n434_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT48), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(new_n704_), .A3(new_n434_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1333gat));
  OR3_X1    g507(.A1(new_n700_), .A2(G71gat), .A3(new_n431_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n696_), .A2(new_n430_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT49), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(G71gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G71gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT109), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n709_), .B(new_n716_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1334gat));
  INV_X1    g517(.A(G78gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n696_), .B2(new_n690_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT50), .Z(new_n721_));
  NAND3_X1  g520(.A1(new_n701_), .A2(new_n719_), .A3(new_n690_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1335gat));
  AND3_X1   g522(.A1(new_n649_), .A2(new_n480_), .A3(new_n695_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n342_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n669_), .A2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n667_), .A2(new_n668_), .A3(KEYINPUT110), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n727_), .A2(new_n480_), .A3(new_n699_), .A4(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n617_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n725_), .B1(new_n730_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g530(.A(G92gat), .B1(new_n724_), .B2(new_n434_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n729_), .A2(new_n403_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G92gat), .ZN(G1337gat));
  NAND4_X1  g533(.A1(new_n649_), .A2(new_n499_), .A3(new_n480_), .A4(new_n695_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(new_n431_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G99gat), .B1(new_n729_), .B2(new_n431_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n738_), .B(new_n739_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1338gat));
  NAND3_X1  g545(.A1(new_n724_), .A2(new_n500_), .A3(new_n692_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n669_), .A2(new_n692_), .A3(new_n480_), .A4(new_n699_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(G106gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G106gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(new_n747_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  INV_X1    g555(.A(KEYINPUT57), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n564_), .B1(new_n558_), .B2(new_n556_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT116), .Z(new_n759_));
  NAND2_X1  g558(.A1(new_n555_), .A2(new_n559_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n565_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n604_), .B2(new_n596_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n579_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n588_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(KEYINPUT55), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT114), .B(new_n768_), .C1(new_n765_), .C2(new_n588_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n586_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n584_), .B1(new_n583_), .B2(new_n571_), .ZN(new_n771_));
  AOI211_X1 g570(.A(KEYINPUT68), .B(KEYINPUT12), .C1(new_n524_), .C2(new_n582_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n580_), .B1(new_n773_), .B2(new_n581_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT114), .B1(new_n774_), .B2(new_n768_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n586_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n766_), .A2(new_n764_), .A3(KEYINPUT55), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n770_), .A2(new_n778_), .A3(new_n598_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(new_n570_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n596_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(KEYINPUT115), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n763_), .B1(new_n781_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n757_), .B1(new_n786_), .B2(new_n613_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n780_), .A2(new_n570_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n779_), .B2(KEYINPUT115), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n782_), .A3(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT57), .B(new_n648_), .C1(new_n790_), .C2(new_n763_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n770_), .A2(new_n778_), .A3(new_n598_), .A4(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n596_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n762_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n796_));
  INV_X1    g595(.A(new_n792_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n779_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n795_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(KEYINPUT118), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(KEYINPUT118), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n794_), .A2(new_n795_), .A3(new_n802_), .A4(new_n798_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n801_), .A2(new_n549_), .A3(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n787_), .A2(new_n791_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n480_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n570_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n479_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n807_), .B2(new_n479_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n653_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT54), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n653_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n806_), .A2(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n434_), .A2(new_n617_), .A3(new_n431_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n393_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(G113gat), .B1(new_n819_), .B2(new_n570_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(KEYINPUT59), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n692_), .B1(new_n806_), .B2(new_n815_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n817_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n821_), .A2(G113gat), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n820_), .B1(new_n825_), .B2(new_n570_), .ZN(G1340gat));
  INV_X1    g625(.A(new_n608_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n821_), .A2(new_n827_), .A3(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT120), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n821_), .A2(new_n830_), .A3(new_n827_), .A4(new_n824_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(G120gat), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n607_), .B2(KEYINPUT60), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT119), .Z(new_n835_));
  OAI211_X1 g634(.A(new_n819_), .B(new_n835_), .C1(KEYINPUT60), .C2(new_n833_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n836_), .ZN(G1341gat));
  AOI21_X1  g636(.A(G127gat), .B1(new_n819_), .B2(new_n479_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n821_), .A2(new_n824_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n479_), .A2(G127gat), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(G1342gat));
  AOI21_X1  g640(.A(G134gat), .B1(new_n819_), .B2(new_n613_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT121), .B(G134gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n653_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n842_), .B1(new_n839_), .B2(new_n844_), .ZN(G1343gat));
  NAND4_X1  g644(.A1(new_n692_), .A2(new_n342_), .A3(new_n403_), .A4(new_n431_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT122), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n806_), .B2(new_n815_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n570_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n827_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n479_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT123), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(KEYINPUT123), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OR3_X1    g657(.A1(new_n855_), .A2(new_n856_), .A3(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1346gat));
  AOI21_X1  g660(.A(G162gat), .B1(new_n848_), .B2(new_n613_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n848_), .A2(new_n549_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(G162gat), .B2(new_n863_), .ZN(G1347gat));
  AND2_X1   g663(.A1(new_n434_), .A2(new_n432_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n570_), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT124), .Z(new_n867_));
  NAND3_X1  g666(.A1(new_n816_), .A2(new_n643_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n868_), .B(G169gat), .C1(KEYINPUT125), .C2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(KEYINPUT125), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n816_), .A2(new_n643_), .A3(new_n865_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n570_), .A3(new_n288_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(G1348gat));
  AND4_X1   g675(.A1(G176gat), .A2(new_n822_), .A3(new_n827_), .A4(new_n865_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n607_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G176gat), .B1(new_n874_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n880_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n877_), .B1(new_n881_), .B2(new_n882_), .ZN(G1349gat));
  NOR3_X1   g682(.A1(new_n873_), .A2(new_n272_), .A3(new_n480_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n822_), .A2(new_n479_), .A3(new_n865_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n266_), .B2(new_n885_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n873_), .B2(new_n653_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n613_), .A2(new_n273_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n873_), .B2(new_n888_), .ZN(G1351gat));
  AOI21_X1  g688(.A(new_n403_), .B1(new_n806_), .B2(new_n815_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n890_), .A2(new_n404_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n570_), .A3(new_n431_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n431_), .A3(new_n827_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g694(.A1(new_n890_), .A2(new_n404_), .A3(new_n431_), .A4(new_n479_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  AND2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n897_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n900_), .A2(KEYINPUT127), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(KEYINPUT127), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n901_), .B2(new_n902_), .ZN(G1354gat));
  AND4_X1   g702(.A1(G218gat), .A2(new_n891_), .A3(new_n431_), .A4(new_n549_), .ZN(new_n904_));
  INV_X1    g703(.A(G218gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n891_), .A2(new_n613_), .A3(new_n431_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1355gat));
endmodule


