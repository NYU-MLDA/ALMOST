//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT34), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT35), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT10), .B(G99gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n209_), .B(new_n210_), .C1(new_n211_), .C2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  OAI22_X1  g012(.A1(KEYINPUT64), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n213_), .A2(new_n214_), .B1(new_n216_), .B2(KEYINPUT9), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT65), .B1(new_n212_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n213_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n209_), .A2(new_n210_), .ZN(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n225_), .A2(KEYINPUT10), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(KEYINPUT10), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n224_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .A4(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(new_n225_), .A3(new_n224_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n232_), .A2(new_n209_), .A3(new_n210_), .A4(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G85gat), .B(G92gat), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT8), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT8), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(new_n238_), .A3(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(G29gat), .A2(G36gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G29gat), .A2(G36gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(G43gat), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G29gat), .ZN(new_n244_));
  INV_X1    g043(.A(G36gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G43gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G29gat), .A2(G36gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n243_), .A2(new_n249_), .A3(G50gat), .ZN(new_n250_));
  INV_X1    g049(.A(G50gat), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n241_), .A2(new_n242_), .A3(G43gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n247_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n230_), .A2(new_n240_), .A3(new_n250_), .A4(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n204_), .A2(new_n205_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT15), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n243_), .A2(new_n249_), .A3(G50gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(G50gat), .B1(new_n243_), .B2(new_n249_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n254_), .A2(KEYINPUT15), .A3(new_n250_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n230_), .A2(new_n240_), .ZN(new_n264_));
  AOI211_X1 g063(.A(new_n206_), .B(new_n257_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n263_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n255_), .A2(KEYINPUT73), .A3(new_n256_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n257_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n265_), .B1(new_n272_), .B2(new_n206_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT74), .B(G134gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G162gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(G190gat), .B(G218gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT36), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT75), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n273_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n277_), .B(KEYINPUT36), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT76), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n273_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(KEYINPUT77), .A2(G22gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(KEYINPUT77), .A2(G22gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G15gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n287_), .A2(G15gat), .A3(new_n288_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G1gat), .B(G8gat), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n291_), .A2(new_n296_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G57gat), .B(G64gat), .Z(new_n301_));
  INV_X1    g100(.A(KEYINPUT11), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G57gat), .B(G64gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n305_));
  XOR2_X1   g104(.A(G71gat), .B(G78gat), .Z(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n305_), .A2(new_n306_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n300_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G231gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n310_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT17), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT16), .B(G183gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(G211gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G155gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  OAI21_X1  g117(.A(new_n313_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(KEYINPUT17), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n319_), .B1(new_n313_), .B2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT78), .Z(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT18), .B(G64gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G92gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G8gat), .B(G36gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT19), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(G169gat), .B2(G176gat), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n334_));
  INV_X1    g133(.A(G169gat), .ZN(new_n335_));
  INV_X1    g134(.A(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G183gat), .ZN(new_n340_));
  INV_X1    g139(.A(G190gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT23), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(G183gat), .A3(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n332_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT92), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G190gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT92), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n348_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n346_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT94), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT83), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n344_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n343_), .A2(KEYINPUT83), .A3(G183gat), .A4(G190gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n342_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(G183gat), .B2(G190gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n335_), .A2(new_n336_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G169gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n365_), .B2(new_n336_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n358_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(new_n358_), .A3(new_n366_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n357_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G211gat), .B(G218gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(G197gat), .B(G204gat), .Z(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(KEYINPUT21), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(KEYINPUT21), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n331_), .B1(new_n370_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n362_), .A2(new_n347_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n355_), .A2(new_n352_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n333_), .A2(new_n337_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT82), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n355_), .A2(new_n352_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n362_), .A2(KEYINPUT84), .A3(new_n347_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n380_), .A2(new_n383_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n366_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n366_), .A2(new_n389_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n345_), .B1(G183gat), .B2(G190gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(new_n375_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n330_), .B1(new_n377_), .B2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n357_), .B(new_n375_), .C1(new_n367_), .C2(new_n369_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n388_), .A2(new_n393_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n376_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n396_), .A2(new_n398_), .A3(KEYINPUT20), .A4(new_n330_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n327_), .B1(new_n395_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n363_), .A2(new_n366_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT94), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n403_), .A2(new_n368_), .B1(new_n346_), .B2(new_n356_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT20), .B(new_n394_), .C1(new_n404_), .C2(new_n375_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n329_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n399_), .A3(new_n326_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n401_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G120gat), .ZN(new_n409_));
  OR2_X1    g208(.A1(G127gat), .A2(G134gat), .ZN(new_n410_));
  INV_X1    g209(.A(G113gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G127gat), .A2(G134gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n411_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n409_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n415_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(G120gat), .A3(new_n413_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT2), .ZN(new_n420_));
  INV_X1    g219(.A(G141gat), .ZN(new_n421_));
  INV_X1    g220(.A(G148gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G155gat), .A2(G162gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT90), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT90), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(new_n433_), .A3(new_n430_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n428_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n430_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n436_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n421_), .A2(new_n422_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n437_), .B(new_n438_), .C1(KEYINPUT1), .C2(new_n431_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n419_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n416_), .A2(new_n418_), .A3(new_n435_), .A4(new_n439_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(KEYINPUT4), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n444_), .B(KEYINPUT95), .Z(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n419_), .A2(new_n446_), .A3(new_n440_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n445_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n441_), .A2(new_n449_), .A3(new_n442_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G1gat), .B(G29gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G57gat), .B(G85gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n448_), .A2(new_n450_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT97), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT97), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n448_), .A2(new_n458_), .A3(new_n450_), .A4(new_n455_), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT98), .B(KEYINPUT33), .Z(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n443_), .A2(new_n449_), .A3(new_n447_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n455_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n441_), .A2(new_n445_), .A3(new_n442_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n456_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n408_), .A2(new_n466_), .A3(KEYINPUT99), .A4(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT99), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n401_), .A2(new_n461_), .A3(new_n407_), .A4(new_n465_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(new_n468_), .ZN(new_n473_));
  OR3_X1    g272(.A1(new_n405_), .A2(KEYINPUT101), .A3(new_n329_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n357_), .A2(KEYINPUT100), .A3(new_n402_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT100), .B1(new_n357_), .B2(new_n402_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n376_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n398_), .A2(KEYINPUT20), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n329_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT101), .B1(new_n405_), .B2(new_n329_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n448_), .A2(new_n450_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n463_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n456_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n406_), .A2(new_n399_), .A3(new_n482_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n484_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n470_), .A2(new_n473_), .A3(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G78gat), .B(G106gat), .Z(new_n491_));
  AND2_X1   g290(.A1(new_n440_), .A2(KEYINPUT29), .ZN(new_n492_));
  INV_X1    g291(.A(G228gat), .ZN(new_n493_));
  INV_X1    g292(.A(G233gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n492_), .A2(new_n375_), .A3(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n495_), .B1(new_n492_), .B2(new_n375_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n491_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n497_), .A3(new_n491_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n440_), .A2(KEYINPUT29), .ZN(new_n502_));
  XOR2_X1   g301(.A(G22gat), .B(G50gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT28), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n502_), .B(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n498_), .B2(KEYINPUT91), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n499_), .A2(KEYINPUT91), .A3(new_n500_), .A4(new_n505_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510_));
  XOR2_X1   g309(.A(G15gat), .B(G43gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(G71gat), .B(G99gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n514_));
  NAND2_X1  g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n513_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n388_), .A2(new_n520_), .A3(new_n393_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n388_), .B2(new_n393_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n519_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n397_), .A2(KEYINPUT30), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(KEYINPUT88), .A3(new_n521_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n518_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT88), .B1(new_n525_), .B2(new_n521_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(new_n517_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n419_), .B(KEYINPUT31), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n527_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n522_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n517_), .B1(new_n533_), .B2(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n524_), .A2(new_n518_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n532_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n510_), .B1(new_n531_), .B2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n530_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n534_), .A2(new_n535_), .A3(new_n532_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(KEYINPUT89), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n490_), .A2(new_n509_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n487_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n407_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n481_), .B2(new_n327_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n401_), .A2(new_n407_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n547_));
  AOI22_X1  g346(.A1(new_n545_), .A2(KEYINPUT27), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n509_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n531_), .A2(new_n536_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n509_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n543_), .B(new_n548_), .C1(new_n549_), .C2(new_n551_), .ZN(new_n552_));
  AOI211_X1 g351(.A(new_n286_), .B(new_n322_), .C1(new_n542_), .C2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT81), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n263_), .A2(KEYINPUT80), .A3(new_n300_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT79), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n254_), .A2(KEYINPUT79), .A3(new_n250_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n560_), .A2(KEYINPUT80), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n263_), .A2(new_n300_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n555_), .B(new_n556_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n555_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n558_), .A2(new_n559_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n300_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n560_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n564_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n335_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(G197gat), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n563_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n563_), .B2(new_n569_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n554_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n572_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n560_), .A2(KEYINPUT80), .B1(new_n263_), .B2(new_n300_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n556_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n564_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n565_), .A2(new_n566_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n555_), .B1(new_n580_), .B2(new_n560_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n576_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n563_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(KEYINPUT81), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n575_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT67), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n309_), .B1(new_n230_), .B2(new_n240_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT68), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n587_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT12), .B1(new_n588_), .B2(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n587_), .B(KEYINPUT12), .C1(new_n588_), .C2(new_n589_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n230_), .A2(new_n240_), .A3(new_n309_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597_));
  INV_X1    g396(.A(G204gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT5), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(G176gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(G176gat), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n588_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT66), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n595_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n593_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n264_), .A2(KEYINPUT66), .A3(new_n308_), .A4(new_n307_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n596_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT69), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n603_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(KEYINPUT69), .A3(new_n601_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n596_), .B2(new_n610_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT13), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n618_), .B1(KEYINPUT70), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n596_), .A2(new_n610_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n616_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n596_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n619_), .A2(KEYINPUT70), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n619_), .A2(KEYINPUT70), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n625_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n586_), .B1(new_n620_), .B2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n553_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n202_), .B1(new_n630_), .B2(new_n487_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT103), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n542_), .A2(new_n552_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT37), .B1(new_n281_), .B2(new_n284_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n273_), .A2(new_n280_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n635_), .B(new_n636_), .C1(new_n273_), .C2(new_n283_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n322_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n633_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n620_), .A2(new_n628_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT71), .Z(new_n642_));
  AND3_X1   g441(.A1(new_n640_), .A2(new_n585_), .A3(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n202_), .A3(new_n487_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT38), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n632_), .A2(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(new_n548_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n553_), .A2(new_n629_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n553_), .A2(KEYINPUT104), .A3(new_n629_), .A4(new_n647_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(G8gat), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n650_), .A2(new_n654_), .A3(G8gat), .A4(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n643_), .A2(new_n292_), .A3(new_n647_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(KEYINPUT40), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  INV_X1    g461(.A(new_n541_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n643_), .A2(new_n290_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n630_), .A2(new_n663_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(new_n665_), .B2(G15gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n664_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT105), .ZN(G1326gat));
  INV_X1    g468(.A(G22gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n509_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n643_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n630_), .A2(new_n671_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G22gat), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT106), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT106), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(KEYINPUT42), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT42), .B1(new_n675_), .B2(new_n676_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n672_), .B1(new_n677_), .B2(new_n678_), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n629_), .A2(new_n322_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n633_), .A2(new_n286_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT110), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n285_), .B1(new_n542_), .B2(new_n552_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(KEYINPUT110), .A3(new_n681_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n244_), .A3(new_n487_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n638_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n542_), .B2(new_n552_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT109), .B1(new_n693_), .B2(KEYINPUT108), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(KEYINPUT109), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n680_), .B(KEYINPUT107), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n692_), .A2(new_n695_), .A3(new_n696_), .A4(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n691_), .B1(new_n633_), .B2(new_n638_), .ZN(new_n699_));
  AOI211_X1 g498(.A(KEYINPUT43), .B(new_n689_), .C1(new_n542_), .C2(new_n552_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n696_), .B(new_n697_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n694_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n543_), .B1(new_n698_), .B2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n688_), .B1(new_n703_), .B2(new_n244_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n684_), .A2(new_n245_), .A3(new_n647_), .A4(new_n686_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT112), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT112), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n709_), .A2(KEYINPUT112), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n709_), .A2(KEYINPUT112), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(KEYINPUT45), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n698_), .A2(new_n702_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n245_), .B1(new_n717_), .B2(new_n647_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n707_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n647_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n721_), .A2(KEYINPUT46), .A3(new_n715_), .A4(new_n712_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1329gat));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n687_), .A2(new_n247_), .A3(new_n663_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n531_), .B(new_n536_), .C1(new_n698_), .C2(new_n702_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n724_), .B(new_n725_), .C1(new_n726_), .C2(new_n247_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n247_), .B1(new_n717_), .B2(new_n550_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n725_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT47), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n727_), .A2(new_n730_), .ZN(G1330gat));
  NAND3_X1  g530(.A1(new_n687_), .A2(new_n251_), .A3(new_n671_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n509_), .B1(new_n698_), .B2(new_n702_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n251_), .ZN(G1331gat));
  NOR2_X1   g533(.A1(new_n641_), .A2(new_n585_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n640_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT113), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n487_), .B1(new_n736_), .B2(KEYINPUT113), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n642_), .A2(new_n585_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n553_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(new_n487_), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n739_), .A2(new_n740_), .B1(new_n743_), .B2(new_n738_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT114), .ZN(G1332gat));
  INV_X1    g544(.A(G64gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n742_), .B2(new_n647_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT48), .Z(new_n748_));
  NAND3_X1  g547(.A1(new_n736_), .A2(new_n746_), .A3(new_n647_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1333gat));
  INV_X1    g549(.A(G71gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n742_), .B2(new_n663_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT49), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n736_), .A2(new_n751_), .A3(new_n663_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1334gat));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n742_), .B2(new_n671_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT50), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n736_), .A2(new_n756_), .A3(new_n671_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1335gat));
  AND3_X1   g559(.A1(new_n741_), .A2(new_n322_), .A3(new_n685_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n487_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n692_), .A2(new_n322_), .A3(new_n735_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(new_n543_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g564(.A(G92gat), .B1(new_n761_), .B2(new_n647_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n647_), .A2(G92gat), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT115), .Z(new_n769_));
  AOI21_X1  g568(.A(new_n766_), .B1(new_n767_), .B2(new_n769_), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n763_), .B2(new_n541_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n761_), .B(new_n550_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g573(.A(G106gat), .B1(new_n763_), .B2(new_n509_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT52), .B(G106gat), .C1(new_n763_), .C2(new_n509_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n761_), .A2(KEYINPUT116), .A3(new_n224_), .A4(new_n671_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n741_), .A2(new_n224_), .A3(new_n322_), .A4(new_n685_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n509_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n777_), .A2(new_n778_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT53), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n777_), .A2(new_n786_), .A3(new_n778_), .A4(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1339gat));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n585_), .B1(new_n620_), .B2(new_n628_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n639_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n639_), .B2(new_n790_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT120), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n564_), .B(new_n556_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n555_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n576_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n796_), .A2(new_n797_), .A3(KEYINPUT118), .A4(new_n576_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n583_), .A3(new_n801_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n618_), .A2(new_n795_), .A3(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n800_), .A2(new_n583_), .A3(new_n801_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT119), .B1(new_n625_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n611_), .B1(new_n575_), .B2(new_n584_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n808_));
  NAND2_X1  g607(.A1(new_n596_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n592_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n608_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n594_), .A2(new_n595_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n812_), .A2(KEYINPUT55), .A3(new_n593_), .A4(new_n592_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n809_), .A2(new_n811_), .A3(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n622_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n814_), .B2(new_n622_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n807_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n286_), .B1(new_n806_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n794_), .B1(new_n818_), .B2(KEYINPUT57), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(KEYINPUT57), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n802_), .A2(new_n611_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT58), .B(new_n821_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n638_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n585_), .A2(new_n624_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n814_), .A2(new_n622_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n622_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n795_), .B1(new_n618_), .B2(new_n802_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n625_), .A2(new_n804_), .A3(KEYINPUT119), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n285_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(KEYINPUT120), .A3(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n819_), .A2(new_n820_), .A3(new_n826_), .A4(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n793_), .B1(new_n839_), .B2(new_n322_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n647_), .A2(new_n543_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n551_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n585_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT59), .B1(new_n840_), .B2(new_n842_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n826_), .B1(new_n837_), .B2(new_n836_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n818_), .A2(KEYINPUT57), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n322_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n791_), .A2(new_n792_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n551_), .A4(new_n841_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n845_), .A2(new_n846_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n846_), .B1(new_n845_), .B2(new_n853_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n586_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n844_), .B1(new_n856_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g656(.A(new_n642_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n845_), .A2(new_n858_), .A3(new_n853_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n843_), .B1(KEYINPUT60), .B2(new_n409_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n409_), .B1(new_n641_), .B2(KEYINPUT60), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT122), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n859_), .A2(new_n409_), .B1(new_n860_), .B2(new_n862_), .ZN(G1341gat));
  INV_X1    g662(.A(new_n322_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G127gat), .B1(new_n843_), .B2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n854_), .A2(new_n855_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n864_), .A2(G127gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(G1342gat));
  AOI21_X1  g667(.A(G134gat), .B1(new_n843_), .B2(new_n286_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n854_), .A2(new_n855_), .A3(new_n689_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g670(.A1(new_n840_), .A2(new_n509_), .A3(new_n663_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n585_), .A3(new_n841_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n858_), .A3(new_n841_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g675(.A1(new_n872_), .A2(new_n864_), .A3(new_n841_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  AND4_X1   g678(.A1(G162gat), .A2(new_n872_), .A3(new_n638_), .A4(new_n841_), .ZN(new_n880_));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n872_), .A2(new_n286_), .A3(new_n841_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n548_), .A2(new_n487_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n663_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n671_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n851_), .A2(new_n886_), .A3(new_n585_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G169gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT123), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n890_), .A3(G169gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n851_), .A2(new_n886_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n851_), .B2(new_n886_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n585_), .B(new_n365_), .C1(new_n897_), .C2(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n889_), .A2(KEYINPUT62), .A3(new_n891_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n894_), .A2(new_n899_), .A3(new_n900_), .ZN(G1348gat));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n851_), .A2(new_n886_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT124), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n641_), .B1(new_n904_), .B2(new_n896_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n902_), .B1(new_n905_), .B2(G176gat), .ZN(new_n906_));
  INV_X1    g705(.A(new_n641_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(KEYINPUT125), .A3(new_n336_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n840_), .A2(new_n671_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n642_), .A2(new_n336_), .A3(new_n885_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n906_), .A2(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(G1349gat));
  AOI21_X1  g711(.A(new_n322_), .B1(new_n904_), .B2(new_n896_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n355_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n910_), .A2(new_n663_), .A3(new_n864_), .A4(new_n884_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n913_), .A2(new_n914_), .B1(new_n915_), .B2(new_n340_), .ZN(G1350gat));
  OAI21_X1  g715(.A(new_n354_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n689_), .B1(new_n904_), .B2(new_n896_), .ZN(new_n918_));
  OAI22_X1  g717(.A1(new_n285_), .A2(new_n917_), .B1(new_n918_), .B2(new_n341_), .ZN(G1351gat));
  NOR2_X1   g718(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT126), .B(G197gat), .Z(new_n921_));
  NAND3_X1  g720(.A1(new_n872_), .A2(new_n585_), .A3(new_n884_), .ZN(new_n922_));
  MUX2_X1   g721(.A(new_n920_), .B(new_n921_), .S(new_n922_), .Z(G1352gat));
  NAND3_X1  g722(.A1(new_n872_), .A2(new_n858_), .A3(new_n884_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g724(.A1(new_n872_), .A2(new_n864_), .A3(new_n884_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  AND2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n926_), .B2(new_n927_), .ZN(G1354gat));
  AND3_X1   g729(.A1(new_n872_), .A2(new_n286_), .A3(new_n884_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n872_), .A2(new_n638_), .A3(new_n884_), .ZN(new_n932_));
  MUX2_X1   g731(.A(new_n931_), .B(new_n932_), .S(G218gat), .Z(G1355gat));
endmodule


