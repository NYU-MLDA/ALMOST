//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT10), .B(G99gat), .Z(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G106gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G85gat), .B(G92gat), .Z(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  OR3_X1    g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT9), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n205_), .A2(new_n208_), .A3(new_n210_), .A4(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n209_), .B1(new_n218_), .B2(new_n204_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n215_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G57gat), .B(G64gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT11), .ZN(new_n224_));
  XOR2_X1   g023(.A(G71gat), .B(G78gat), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n223_), .A2(KEYINPUT11), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n224_), .A2(new_n225_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n214_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n230_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT12), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT68), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n241_), .A3(new_n238_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n233_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n222_), .A2(KEYINPUT66), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n236_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n230_), .A2(KEYINPUT12), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n244_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT67), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n244_), .A2(new_n246_), .A3(new_n251_), .A4(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G230gat), .A2(G233gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n243_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n232_), .A2(KEYINPUT65), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n237_), .B1(new_n232_), .B2(KEYINPUT65), .ZN(new_n257_));
  OAI211_X1 g056(.A(G230gat), .B(G233gat), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G120gat), .B(G148gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT5), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G176gat), .B(G204gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n255_), .A2(new_n258_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT69), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n255_), .A2(new_n266_), .A3(new_n258_), .A4(new_n263_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n255_), .A2(new_n258_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n262_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT13), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n268_), .A2(KEYINPUT13), .A3(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT70), .ZN(new_n276_));
  XOR2_X1   g075(.A(G78gat), .B(G106gat), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G141gat), .A2(G148gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT2), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n283_), .A2(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT91), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT91), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n291_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT92), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n281_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n288_), .A2(new_n293_), .A3(KEYINPUT92), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n280_), .A2(KEYINPUT1), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(G155gat), .A3(G162gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n300_), .A3(new_n279_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G141gat), .B(G148gat), .Z(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT90), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n301_), .A2(new_n302_), .A3(KEYINPUT90), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n296_), .A2(new_n297_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G211gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(G218gat), .ZN(new_n311_));
  INV_X1    g110(.A(G218gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n312_), .A2(G211gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT95), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(G211gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(G218gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT95), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G197gat), .A2(G204gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT21), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n314_), .A2(new_n318_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT96), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n314_), .A2(new_n322_), .A3(KEYINPUT96), .A4(new_n318_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n314_), .A2(new_n318_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n322_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(KEYINPUT93), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT93), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT21), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n333_), .A2(new_n334_), .A3(KEYINPUT94), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT94), .B1(new_n333_), .B2(new_n334_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n328_), .B(new_n329_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n327_), .A2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(G228gat), .B(G233gat), .C1(new_n309_), .C2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n294_), .A2(new_n295_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n281_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n297_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n305_), .A2(new_n306_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT29), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n317_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT96), .B1(new_n348_), .B2(new_n322_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n326_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n337_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT97), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT97), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n327_), .A2(new_n353_), .A3(new_n337_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G228gat), .A2(G233gat), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n345_), .A2(new_n352_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n278_), .B1(new_n339_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n307_), .A2(new_n360_), .A3(new_n308_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n359_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT28), .B1(new_n344_), .B2(KEYINPUT29), .ZN(new_n365_));
  INV_X1    g164(.A(new_n359_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n339_), .A2(new_n278_), .A3(new_n356_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n358_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n367_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n339_), .A2(new_n278_), .A3(new_n356_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(new_n357_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT18), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380_));
  OR3_X1    g179(.A1(new_n380_), .A2(KEYINPUT82), .A3(G169gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT84), .B(G176gat), .ZN(new_n382_));
  INV_X1    g181(.A(G169gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT22), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT82), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n381_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n380_), .A2(G169gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT83), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n386_), .A2(new_n388_), .B1(G169gat), .B2(G176gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT23), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(G183gat), .B2(G190gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n389_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT26), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G190gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT25), .B(G183gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT26), .B(G190gat), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n403_), .B(new_n404_), .C1(new_n405_), .C2(new_n402_), .ZN(new_n406_));
  OR2_X1    g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(KEYINPUT24), .A3(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n407_), .A2(KEYINPUT24), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n406_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT23), .B1(new_n393_), .B2(new_n394_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n390_), .B1(G183gat), .B2(G190gat), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n399_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n352_), .A2(new_n354_), .A3(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT20), .ZN(new_n422_));
  INV_X1    g221(.A(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT26), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n401_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G183gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT25), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT25), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G183gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n409_), .B1(new_n425_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT99), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n395_), .A2(new_n410_), .A3(new_n396_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT99), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n434_), .B(new_n409_), .C1(new_n425_), .C2(new_n430_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n432_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  OAI22_X1  g235(.A1(new_n413_), .A2(new_n414_), .B1(G183gat), .B2(G190gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT100), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n387_), .A2(new_n384_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n387_), .B2(new_n384_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n382_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n441_), .A3(new_n408_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n327_), .A2(new_n436_), .A3(new_n337_), .A4(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT101), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n422_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n436_), .A2(new_n442_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n338_), .A2(new_n446_), .A3(KEYINPUT101), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n418_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n398_), .A2(new_n389_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n327_), .A2(new_n353_), .A3(new_n337_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n353_), .B1(new_n327_), .B2(new_n337_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n436_), .A2(new_n442_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n351_), .B2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n421_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n379_), .B1(new_n448_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT102), .ZN(new_n458_));
  INV_X1    g257(.A(new_n421_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n417_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n455_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n418_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n378_), .A3(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n457_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  OAI211_X1 g265(.A(KEYINPUT102), .B(new_n379_), .C1(new_n448_), .C2(new_n456_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n453_), .B1(new_n338_), .B2(new_n446_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n418_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n459_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n452_), .A2(new_n455_), .A3(new_n421_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(KEYINPUT27), .B(new_n464_), .C1(new_n473_), .C2(new_n378_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n374_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G127gat), .B(G134gat), .Z(new_n476_));
  XOR2_X1   g275(.A(G113gat), .B(G120gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT30), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n417_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n449_), .A2(KEYINPUT30), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G71gat), .B(G99gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT85), .B(G43gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n485_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G227gat), .ZN(new_n490_));
  INV_X1    g289(.A(G233gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n487_), .B(new_n488_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT86), .B(G15gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n493_), .A2(new_n496_), .A3(new_n494_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n482_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n480_), .A2(new_n481_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n500_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n496_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT87), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT31), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n503_), .A2(new_n508_), .A3(new_n509_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT88), .B1(new_n482_), .B2(new_n502_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n513_), .B2(new_n508_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n478_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n478_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n344_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n307_), .A2(new_n478_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT4), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G225gat), .A2(G233gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR4_X1   g320(.A1(new_n307_), .A2(KEYINPUT103), .A3(KEYINPUT4), .A4(new_n478_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT103), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n478_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n519_), .B(new_n521_), .C1(new_n522_), .C2(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n342_), .A2(new_n343_), .A3(new_n478_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n520_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G1gat), .B(G29gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G85gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT104), .B(KEYINPUT0), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n529_), .B2(new_n520_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n531_), .A2(new_n537_), .B1(new_n527_), .B2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n504_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n509_), .B1(new_n504_), .B2(new_n501_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT31), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(new_n511_), .A3(new_n516_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n515_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n475_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n370_), .A2(new_n373_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n468_), .A2(new_n539_), .A3(new_n546_), .A4(new_n474_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n465_), .A2(new_n467_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n517_), .A2(new_n518_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n537_), .B1(new_n549_), .B2(new_n520_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n522_), .A2(new_n526_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n521_), .B1(new_n529_), .B2(KEYINPUT4), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n527_), .A2(new_n538_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT33), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT33), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n527_), .A2(new_n556_), .A3(new_n538_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n553_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n531_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n554_), .B1(new_n559_), .B2(new_n536_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n378_), .A2(KEYINPUT32), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n462_), .A2(new_n463_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n548_), .A2(new_n558_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n547_), .B1(new_n565_), .B2(new_n546_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n542_), .A2(new_n511_), .A3(new_n516_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n516_), .B1(new_n542_), .B2(new_n511_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n515_), .A2(KEYINPUT89), .A3(new_n543_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n545_), .B1(new_n566_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G1gat), .ZN(new_n574_));
  INV_X1    g373(.A(G8gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n577_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G15gat), .B(G22gat), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G1gat), .B(G8gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT77), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n583_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G29gat), .B(G36gat), .Z(new_n587_));
  XOR2_X1   g386(.A(G43gat), .B(G50gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n586_), .B(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n586_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n589_), .B(KEYINPUT15), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n586_), .A2(new_n589_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n591_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n593_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n573_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT78), .Z(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n586_), .A2(new_n230_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n586_), .A2(new_n230_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT16), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT17), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n614_), .A2(new_n616_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT79), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n614_), .A2(new_n616_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT17), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n620_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n624_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n244_), .A2(new_n246_), .A3(new_n595_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT35), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT34), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n222_), .A2(new_n589_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n636_), .A2(new_n633_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n632_), .B(new_n637_), .C1(new_n633_), .C2(new_n636_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT71), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT36), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT74), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n642_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT73), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT37), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT75), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n646_), .A2(KEYINPUT36), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT72), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n640_), .A2(new_n641_), .A3(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n649_), .A2(new_n653_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n653_), .B1(new_n649_), .B2(new_n656_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n652_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n649_), .A2(new_n656_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT75), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n662_), .A2(KEYINPUT37), .A3(new_n651_), .A4(new_n657_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n631_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n276_), .A2(new_n607_), .A3(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n574_), .A3(new_n560_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n606_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n661_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n573_), .A2(new_n670_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n268_), .A2(KEYINPUT13), .A3(new_n270_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT13), .B1(new_n268_), .B2(new_n270_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n622_), .A2(new_n623_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n630_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(new_n625_), .ZN(new_n677_));
  AND4_X1   g476(.A1(new_n669_), .A2(new_n671_), .A3(new_n674_), .A4(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n574_), .B1(new_n678_), .B2(new_n560_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n668_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n680_), .B1(new_n667_), .B2(new_n666_), .ZN(G1324gat));
  NAND2_X1  g480(.A1(new_n468_), .A2(new_n474_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n575_), .B1(new_n678_), .B2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT39), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n665_), .A2(new_n575_), .A3(new_n682_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g486(.A(G15gat), .ZN(new_n688_));
  INV_X1    g487(.A(new_n572_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n678_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT41), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n665_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1326gat));
  INV_X1    g492(.A(G22gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n678_), .B2(new_n546_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n546_), .A2(new_n694_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT106), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n665_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1327gat));
  AOI21_X1  g500(.A(KEYINPUT110), .B1(new_n670_), .B2(new_n631_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n677_), .A2(new_n661_), .A3(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n672_), .A2(new_n705_), .A3(new_n673_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n607_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G29gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n560_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n273_), .A2(new_n669_), .A3(new_n274_), .A4(new_n631_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n566_), .A2(new_n572_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n545_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n660_), .A2(new_n663_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n713_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(KEYINPUT107), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n573_), .A2(new_n717_), .A3(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n712_), .C1(new_n719_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n721_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n716_), .A2(new_n718_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n713_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(new_n573_), .B2(new_n717_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n711_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n727_), .A2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n712_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n725_), .A2(new_n731_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n560_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n710_), .B1(new_n736_), .B2(G29gat), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT109), .B(new_n708_), .C1(new_n735_), .C2(new_n560_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n709_), .B1(new_n737_), .B2(new_n738_), .ZN(G1328gat));
  INV_X1    g538(.A(KEYINPUT116), .ZN(new_n740_));
  INV_X1    g539(.A(G36gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n725_), .A2(new_n731_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n682_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n734_), .B2(new_n732_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n741_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n745_));
  XOR2_X1   g544(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n746_));
  NOR2_X1   g545(.A1(new_n743_), .A2(G36gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n607_), .A2(new_n706_), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n607_), .A2(new_n706_), .A3(KEYINPUT112), .A4(new_n747_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n746_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n746_), .A3(new_n751_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT113), .B1(new_n745_), .B2(new_n755_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n750_), .A2(new_n746_), .A3(new_n751_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(new_n752_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n682_), .B1(new_n730_), .B2(KEYINPUT44), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n725_), .B2(new_n731_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n758_), .B(new_n759_), .C1(new_n761_), .C2(new_n741_), .ZN(new_n762_));
  XOR2_X1   g561(.A(KEYINPUT114), .B(KEYINPUT46), .Z(new_n763_));
  AND3_X1   g562(.A1(new_n756_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n758_), .B(KEYINPUT46), .C1(new_n761_), .C2(new_n741_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n723_), .A2(new_n724_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT108), .B1(new_n730_), .B2(KEYINPUT44), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n744_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(G36gat), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n771_), .A2(KEYINPUT115), .A3(KEYINPUT46), .A4(new_n758_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n767_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n740_), .B1(new_n764_), .B2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n756_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n775_), .A2(KEYINPUT116), .A3(new_n767_), .A4(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1329gat));
  NOR2_X1   g576(.A1(new_n568_), .A2(new_n569_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n735_), .A2(G43gat), .A3(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n707_), .A2(new_n689_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(G43gat), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(KEYINPUT117), .B(KEYINPUT47), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(G1330gat));
  AOI21_X1  g582(.A(G50gat), .B1(new_n707_), .B2(new_n546_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n546_), .A2(G50gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n735_), .B2(new_n785_), .ZN(G1331gat));
  INV_X1    g585(.A(G57gat), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n276_), .A2(new_n669_), .A3(new_n631_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(new_n671_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n789_), .B2(new_n560_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n716_), .A2(new_n275_), .A3(new_n606_), .A4(new_n664_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT118), .Z(new_n792_));
  AND3_X1   g591(.A1(new_n792_), .A2(new_n787_), .A3(new_n560_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1332gat));
  INV_X1    g593(.A(G64gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n789_), .B2(new_n682_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT48), .Z(new_n797_));
  NAND3_X1  g596(.A1(new_n792_), .A2(new_n795_), .A3(new_n682_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1333gat));
  INV_X1    g598(.A(G71gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n789_), .B2(new_n689_), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT49), .Z(new_n802_));
  NAND3_X1  g601(.A1(new_n792_), .A2(new_n800_), .A3(new_n689_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1334gat));
  INV_X1    g603(.A(G78gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n789_), .B2(new_n546_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT50), .Z(new_n807_));
  NAND3_X1  g606(.A1(new_n792_), .A2(new_n805_), .A3(new_n546_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1335gat));
  NOR4_X1   g608(.A1(new_n276_), .A2(new_n573_), .A3(new_n669_), .A4(new_n705_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n211_), .A3(new_n560_), .ZN(new_n811_));
  AND4_X1   g610(.A1(new_n606_), .A2(new_n733_), .A3(new_n275_), .A4(new_n631_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(new_n560_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n813_), .B2(new_n211_), .ZN(G1336gat));
  NAND3_X1  g613(.A1(new_n810_), .A2(new_n212_), .A3(new_n682_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n812_), .A2(new_n682_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(new_n212_), .ZN(G1337gat));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n689_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n778_), .A2(new_n206_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n818_), .A2(G99gat), .B1(new_n810_), .B2(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT119), .B(KEYINPUT51), .Z(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n823_), .B(new_n824_), .C1(new_n825_), .C2(new_n820_), .ZN(G1338gat));
  INV_X1    g625(.A(G106gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n812_), .B2(new_n546_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n810_), .A2(new_n546_), .A3(new_n207_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g632(.A1(new_n590_), .A2(new_n591_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n596_), .A2(new_n597_), .A3(new_n592_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n603_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n605_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n254_), .B1(new_n243_), .B2(new_n253_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n255_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n243_), .A2(new_n253_), .A3(KEYINPUT55), .A4(new_n254_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(KEYINPUT56), .A3(new_n262_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT56), .B1(new_n843_), .B2(new_n262_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n268_), .B(new_n838_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n717_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n268_), .A2(new_n669_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n846_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n844_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n837_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n661_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n849_), .A2(new_n850_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n855_), .A2(new_n856_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n669_), .B(new_n631_), .C1(new_n660_), .C2(new_n663_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n674_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n674_), .A2(new_n606_), .A3(new_n664_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(KEYINPUT54), .ZN(new_n867_));
  AOI211_X1 g666(.A(KEYINPUT122), .B(new_n861_), .C1(new_n860_), .C2(new_n674_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n859_), .A2(new_n631_), .B1(new_n864_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n475_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n560_), .A3(new_n778_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(G113gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n669_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n872_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n864_), .A2(new_n869_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n677_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT59), .B(new_n878_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n606_), .B1(new_n877_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n875_), .B1(new_n882_), .B2(new_n874_), .ZN(G1340gat));
  INV_X1    g682(.A(G120gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n674_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n873_), .B(new_n885_), .C1(KEYINPUT60), .C2(new_n884_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n276_), .B1(new_n877_), .B2(new_n881_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G120gat), .B1(new_n887_), .B2(new_n888_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n886_), .B1(new_n889_), .B2(new_n890_), .ZN(G1341gat));
  NOR3_X1   g690(.A1(new_n870_), .A2(new_n631_), .A3(new_n872_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n892_), .A2(new_n893_), .A3(G127gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n892_), .B2(G127gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n877_), .A2(new_n881_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n677_), .A2(G127gat), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n894_), .A2(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1342gat));
  INV_X1    g697(.A(G134gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n873_), .A2(new_n899_), .A3(new_n670_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n717_), .B1(new_n877_), .B2(new_n881_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1343gat));
  INV_X1    g701(.A(new_n870_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n689_), .A2(new_n539_), .A3(new_n374_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(new_n743_), .A3(new_n904_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n905_), .A2(new_n606_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G141gat), .ZN(G1344gat));
  OR2_X1    g706(.A1(new_n905_), .A2(new_n276_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g708(.A1(new_n905_), .A2(new_n631_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT61), .B(G155gat), .Z(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1346gat));
  OAI21_X1  g711(.A(G162gat), .B1(new_n905_), .B2(new_n717_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n661_), .A2(G162gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n905_), .B2(new_n914_), .ZN(G1347gat));
  NOR4_X1   g714(.A1(new_n572_), .A2(new_n560_), .A3(new_n743_), .A4(new_n546_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n903_), .A2(new_n669_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n917_), .A2(new_n918_), .A3(G169gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n903_), .A2(new_n916_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n921_), .B(new_n669_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n918_), .B1(new_n917_), .B2(G169gat), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n919_), .B1(new_n922_), .B2(new_n923_), .ZN(G1348gat));
  INV_X1    g723(.A(new_n276_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(G176gat), .ZN(new_n926_));
  OR3_X1    g725(.A1(new_n920_), .A2(KEYINPUT125), .A3(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT125), .B1(new_n920_), .B2(new_n926_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n921_), .A2(new_n275_), .ZN(new_n929_));
  AOI22_X1  g728(.A1(new_n927_), .A2(new_n928_), .B1(new_n929_), .B2(new_n382_), .ZN(G1349gat));
  NOR2_X1   g729(.A1(new_n920_), .A2(new_n631_), .ZN(new_n931_));
  MUX2_X1   g730(.A(G183gat), .B(new_n404_), .S(new_n931_), .Z(G1350gat));
  NAND3_X1  g731(.A1(new_n921_), .A2(new_n405_), .A3(new_n670_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n903_), .A2(new_n718_), .A3(new_n916_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n934_), .A2(new_n935_), .A3(G190gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n934_), .B2(G190gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n933_), .B1(new_n936_), .B2(new_n937_), .ZN(G1351gat));
  NOR2_X1   g737(.A1(new_n374_), .A2(new_n560_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n572_), .A2(new_n939_), .A3(new_n682_), .ZN(new_n940_));
  OAI21_X1  g739(.A(KEYINPUT127), .B1(new_n870_), .B2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942_));
  INV_X1    g741(.A(new_n940_), .ZN(new_n943_));
  OAI211_X1 g742(.A(new_n942_), .B(new_n943_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n941_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n669_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n925_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  AND4_X1   g750(.A1(new_n677_), .A2(new_n945_), .A3(new_n950_), .A4(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n950_), .B1(new_n945_), .B2(new_n677_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1354gat));
  NAND3_X1  g753(.A1(new_n945_), .A2(new_n312_), .A3(new_n670_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n717_), .B1(new_n941_), .B2(new_n944_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n312_), .ZN(G1355gat));
endmodule


