//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_;
  INV_X1    g000(.A(G230gat), .ZN(new_n202_));
  INV_X1    g001(.A(G233gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n205_));
  NOR2_X1   g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  INV_X1    g006(.A(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(G92gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n205_), .A2(new_n207_), .A3(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n205_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT10), .B(G99gat), .Z(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT6), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n211_), .A2(new_n212_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT66), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT7), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n223_), .A2(new_n219_), .A3(new_n220_), .A4(KEYINPUT66), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n217_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(KEYINPUT67), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n210_), .A2(new_n206_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n225_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n218_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G78gat), .Z(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n235_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n218_), .B(new_n239_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(KEYINPUT12), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT12), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n232_), .A2(new_n244_), .A3(new_n240_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n204_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n242_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n204_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G120gat), .B(G148gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G176gat), .B(G204gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n255_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n247_), .A2(new_n249_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n260_));
  NAND2_X1  g059(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(new_n258_), .A3(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G29gat), .B(G36gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G43gat), .B(G50gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT15), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n232_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G232gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT35), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n268_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n270_), .B(new_n275_), .C1(new_n232_), .C2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n273_), .A2(new_n274_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G190gat), .B(G218gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G134gat), .B(G162gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(KEYINPUT36), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n278_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n279_), .A2(new_n284_), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n282_), .B(KEYINPUT36), .Z(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT37), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n287_), .A2(KEYINPUT37), .A3(new_n290_), .ZN(new_n294_));
  AND2_X1   g093(.A1(G231gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n239_), .B(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G15gat), .B(G22gat), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G8gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT72), .B(G1gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n300_), .A2(G8gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT14), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n298_), .B(new_n299_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n299_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n302_), .B1(new_n300_), .B2(G8gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(new_n297_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n296_), .B(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G127gat), .B(G155gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT16), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G183gat), .B(G211gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT17), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n312_), .A2(new_n313_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n308_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT73), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n315_), .B(new_n320_), .C1(new_n317_), .C2(new_n308_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n319_), .A2(new_n321_), .A3(KEYINPUT74), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT74), .B1(new_n319_), .B2(new_n321_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AND4_X1   g123(.A1(new_n265_), .A2(new_n293_), .A3(new_n294_), .A4(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n325_), .B(KEYINPUT75), .Z(new_n326_));
  NOR2_X1   g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n328_), .B2(KEYINPUT1), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT90), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G141gat), .A3(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n329_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT91), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n329_), .A2(new_n334_), .A3(KEYINPUT91), .A4(new_n337_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n332_), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n330_), .A2(KEYINPUT90), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n343_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT92), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n346_), .A2(new_n351_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n335_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(new_n328_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n342_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT28), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n340_), .A2(new_n341_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n360_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G22gat), .B(G50gat), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n360_), .B1(new_n342_), .B2(new_n359_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(KEYINPUT21), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT21), .ZN(new_n377_));
  AND2_X1   g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(new_n373_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G211gat), .B(G218gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n378_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G211gat), .B(G218gat), .Z(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n381_), .A2(new_n384_), .A3(KEYINPUT93), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT93), .B1(new_n381_), .B2(new_n384_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n371_), .B1(new_n372_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n381_), .A2(new_n384_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n370_), .B(new_n391_), .C1(new_n363_), .C2(new_n360_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n392_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n389_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n369_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(KEYINPUT94), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT94), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n388_), .A2(new_n398_), .A3(new_n390_), .A4(new_n392_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n369_), .A2(new_n397_), .A3(new_n395_), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT95), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n390_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n403_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n404_), .A2(KEYINPUT95), .A3(new_n399_), .A4(new_n397_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n396_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(KEYINPUT19), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT96), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT81), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(G169gat), .A3(G176gat), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n412_), .A2(new_n414_), .A3(KEYINPUT24), .ZN(new_n415_));
  INV_X1    g214(.A(G169gat), .ZN(new_n416_));
  INV_X1    g215(.A(G176gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(KEYINPUT80), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(G169gat), .B2(G176gat), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n415_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G183gat), .ZN(new_n424_));
  INV_X1    g223(.A(G190gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT23), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n424_), .A2(KEYINPUT23), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(G190gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT23), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n427_), .A2(new_n430_), .A3(G183gat), .A4(G190gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n426_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n418_), .A2(new_n420_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT24), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT26), .B(G190gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT25), .B(G183gat), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n434_), .A2(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n412_), .A2(new_n414_), .A3(KEYINPUT24), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT82), .B1(new_n439_), .B2(new_n434_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n423_), .A2(new_n433_), .A3(new_n438_), .A4(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n412_), .A2(new_n414_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n430_), .A2(G183gat), .A3(G190gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n426_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G183gat), .A2(G190gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT22), .B(G169gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT84), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n449_), .B1(new_n416_), .B2(KEYINPUT22), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n417_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n447_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n441_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT20), .B1(new_n454_), .B2(new_n391_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n391_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n433_), .A2(KEYINPUT99), .A3(new_n446_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT99), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n430_), .B1(G183gat), .B2(G190gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n443_), .A2(KEYINPUT83), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(new_n431_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n458_), .B1(new_n461_), .B2(new_n445_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n442_), .B1(new_n417_), .B2(new_n448_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n411_), .A2(KEYINPUT24), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n465_), .A2(KEYINPUT98), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(KEYINPUT98), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n421_), .A3(new_n467_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n434_), .A2(new_n435_), .B1(new_n426_), .B2(new_n443_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n437_), .B(KEYINPUT97), .ZN(new_n470_));
  INV_X1    g269(.A(new_n436_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n468_), .B(new_n469_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n456_), .B1(new_n464_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n410_), .B1(new_n455_), .B2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G8gat), .B(G36gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n454_), .B2(new_n391_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n464_), .A2(new_n456_), .A3(new_n472_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n409_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n474_), .A2(new_n479_), .A3(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n484_), .A2(KEYINPUT27), .ZN(new_n485_));
  INV_X1    g284(.A(new_n479_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n455_), .A2(new_n473_), .A3(new_n410_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n387_), .A2(new_n464_), .A3(new_n472_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n409_), .B1(new_n481_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT104), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(KEYINPUT104), .B(new_n486_), .C1(new_n487_), .C2(new_n489_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT27), .ZN(new_n495_));
  INV_X1    g294(.A(new_n484_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n479_), .B1(new_n474_), .B2(new_n483_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n407_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G127gat), .B(G134gat), .Z(new_n501_));
  XOR2_X1   g300(.A(G113gat), .B(G120gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT31), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT86), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n441_), .A2(KEYINPUT30), .A3(new_n453_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT30), .B1(new_n441_), .B2(new_n453_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n505_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(KEYINPUT86), .A3(new_n506_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G227gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT85), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G71gat), .B(G99gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G15gat), .B(G43gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n509_), .A2(new_n511_), .A3(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n510_), .A2(new_n517_), .A3(KEYINPUT86), .A4(new_n506_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT87), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n504_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n504_), .A2(new_n522_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n519_), .B(new_n520_), .C1(KEYINPUT87), .C2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n342_), .A2(new_n359_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n503_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n363_), .A2(new_n503_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G225gat), .A2(G233gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n531_), .B(KEYINPUT101), .Z(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G1gat), .B(G29gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G57gat), .B(G85gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n342_), .A2(new_n359_), .A3(new_n503_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n503_), .B1(new_n342_), .B2(new_n359_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT4), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n527_), .A2(new_n542_), .A3(new_n528_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n532_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n534_), .B(new_n539_), .C1(new_n543_), .C2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n529_), .A2(new_n530_), .A3(KEYINPUT4), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n533_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n539_), .B1(new_n550_), .B2(new_n534_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n526_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n500_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n523_), .A2(new_n557_), .A3(new_n525_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n479_), .A2(KEYINPUT32), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n474_), .A2(new_n561_), .A3(new_n483_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n562_), .B(new_n564_), .C1(new_n547_), .C2(new_n551_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT103), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n544_), .A2(new_n533_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n543_), .B2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n540_), .A2(new_n541_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n539_), .B1(new_n569_), .B2(new_n532_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n548_), .A2(KEYINPUT103), .A3(new_n533_), .A4(new_n544_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n568_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n546_), .A2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n550_), .A2(KEYINPUT33), .A3(new_n534_), .A4(new_n539_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n497_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n484_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n565_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n406_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n494_), .A2(new_n552_), .A3(new_n498_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n406_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n560_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT105), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n406_), .A2(new_n579_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n406_), .B2(new_n581_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT105), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n560_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n556_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G169gat), .B(G197gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n307_), .A2(new_n268_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT76), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G229gat), .A2(G233gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n269_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n276_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n594_), .A2(KEYINPUT76), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT76), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n307_), .B2(new_n268_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n599_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT77), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT77), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n599_), .B(new_n605_), .C1(new_n600_), .C2(new_n602_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n596_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT78), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n598_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  AOI211_X1 g408(.A(KEYINPUT78), .B(new_n596_), .C1(new_n604_), .C2(new_n606_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n593_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n596_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n605_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n606_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n612_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT78), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n607_), .A2(new_n608_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n616_), .A2(new_n617_), .A3(new_n598_), .A4(new_n592_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n618_), .A3(KEYINPUT79), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT79), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n620_), .B(new_n593_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n589_), .A2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n326_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n552_), .A2(new_n300_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT38), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n291_), .B(KEYINPUT107), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n589_), .A2(KEYINPUT108), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT108), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n586_), .A2(new_n587_), .A3(new_n560_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n587_), .B1(new_n586_), .B2(new_n560_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n555_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n631_), .B1(new_n634_), .B2(new_n628_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n630_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n265_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n319_), .A2(new_n321_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n637_), .A2(new_n622_), .A3(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT106), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(new_n553_), .ZN(new_n642_));
  INV_X1    g441(.A(G1gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n627_), .B1(new_n642_), .B2(new_n643_), .ZN(G1324gat));
  INV_X1    g443(.A(G8gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n624_), .A2(new_n645_), .A3(new_n499_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n640_), .B(new_n499_), .C1(new_n630_), .C2(new_n635_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(new_n648_), .A3(G8gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G8gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n646_), .B(new_n652_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  INV_X1    g455(.A(G15gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n560_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n624_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n640_), .B(new_n658_), .C1(new_n630_), .C2(new_n635_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT41), .B1(new_n660_), .B2(G15gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT110), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT110), .B(new_n659_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1326gat));
  INV_X1    g466(.A(G22gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n624_), .A2(new_n668_), .A3(new_n407_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n641_), .A2(new_n407_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(G22gat), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT42), .B(new_n668_), .C1(new_n641_), .C2(new_n407_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(G1327gat));
  NOR3_X1   g473(.A1(new_n637_), .A2(new_n291_), .A3(new_n324_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n623_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n553_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n637_), .A2(new_n622_), .A3(new_n324_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n293_), .A2(new_n294_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n589_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n634_), .B2(new_n679_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n678_), .B1(new_n682_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT44), .B(new_n678_), .C1(new_n682_), .C2(new_n685_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n553_), .A2(G29gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n677_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n499_), .A3(new_n689_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(new_n622_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n499_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(G36gat), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n634_), .A2(new_n699_), .A3(new_n675_), .A4(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT45), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT45), .ZN(new_n704_));
  OAI22_X1  g503(.A1(new_n703_), .A2(new_n704_), .B1(KEYINPUT112), .B2(KEYINPUT46), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n696_), .B1(new_n698_), .B2(new_n706_), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n695_), .B(new_n705_), .C1(new_n697_), .C2(G36gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(G43gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n526_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n688_), .A2(new_n689_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n676_), .A2(new_n658_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g515(.A(G50gat), .B1(new_n676_), .B2(new_n407_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n407_), .A2(G50gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n690_), .B2(new_n718_), .ZN(G1331gat));
  INV_X1    g518(.A(G57gat), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n637_), .A2(new_n622_), .A3(new_n324_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n636_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(new_n553_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n680_), .A2(new_n324_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n637_), .A2(new_n622_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n589_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(new_n720_), .A3(new_n553_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n723_), .A2(new_n727_), .ZN(G1332gat));
  INV_X1    g527(.A(G64gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n729_), .A3(new_n499_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n722_), .A2(new_n499_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(G64gat), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT48), .B(new_n729_), .C1(new_n722_), .C2(new_n499_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(G1333gat));
  NOR2_X1   g534(.A1(new_n560_), .A2(G71gat), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT114), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n726_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n722_), .A2(new_n658_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(G71gat), .ZN(new_n741_));
  INV_X1    g540(.A(G71gat), .ZN(new_n742_));
  INV_X1    g541(.A(new_n739_), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n742_), .B(new_n743_), .C1(new_n722_), .C2(new_n658_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n738_), .B1(new_n741_), .B2(new_n744_), .ZN(G1334gat));
  INV_X1    g544(.A(G78gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n726_), .A2(new_n746_), .A3(new_n407_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n722_), .A2(new_n407_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(G78gat), .ZN(new_n750_));
  INV_X1    g549(.A(new_n748_), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n746_), .B(new_n751_), .C1(new_n722_), .C2(new_n407_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n750_), .B2(new_n752_), .ZN(G1335gat));
  NOR4_X1   g552(.A1(new_n589_), .A2(new_n291_), .A3(new_n324_), .A4(new_n725_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n553_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n208_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n756_), .A2(KEYINPUT116), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(KEYINPUT116), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n682_), .A2(new_n685_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n699_), .A2(new_n265_), .A3(new_n324_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n552_), .A2(new_n208_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT117), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n757_), .A2(new_n758_), .B1(new_n761_), .B2(new_n763_), .ZN(G1336gat));
  NAND3_X1  g563(.A1(new_n754_), .A2(new_n209_), .A3(new_n499_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n761_), .A2(new_n499_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n209_), .ZN(G1337gat));
  NAND4_X1  g566(.A1(new_n754_), .A2(new_n213_), .A3(new_n525_), .A4(new_n523_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n759_), .A2(new_n658_), .A3(new_n760_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n219_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT51), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n768_), .C1(new_n769_), .C2(new_n219_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n754_), .A2(new_n214_), .A3(new_n407_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n407_), .B(new_n760_), .C1(new_n682_), .C2(new_n685_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G106gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G106gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n775_), .B(new_n781_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1339gat));
  XNOR2_X1  g584(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n325_), .A2(new_n622_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT120), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT120), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n325_), .A2(new_n789_), .A3(new_n622_), .A4(new_n786_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n325_), .A2(new_n622_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n788_), .B(new_n790_), .C1(new_n791_), .C2(new_n786_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n612_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n593_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT121), .B1(new_n793_), .B2(new_n592_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n595_), .A2(new_n612_), .A3(new_n597_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n799_), .A2(new_n618_), .A3(new_n258_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n243_), .A2(new_n204_), .A3(new_n245_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n247_), .A2(KEYINPUT55), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n257_), .B1(new_n246_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT122), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n802_), .A2(new_n804_), .A3(KEYINPUT122), .A4(KEYINPUT56), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  INV_X1    g608(.A(new_n801_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n810_), .A2(new_n246_), .A3(new_n803_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n246_), .A2(new_n803_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n255_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n807_), .A2(new_n808_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n800_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n800_), .A2(KEYINPUT58), .A3(new_n815_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n679_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  INV_X1    g620(.A(new_n258_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n814_), .B2(new_n805_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n619_), .A2(new_n621_), .A3(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n799_), .A2(new_n618_), .A3(new_n259_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n821_), .B1(new_n826_), .B2(new_n291_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n291_), .ZN(new_n828_));
  AOI211_X1 g627(.A(KEYINPUT57), .B(new_n828_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n820_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n792_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n526_), .A2(new_n552_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n500_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(new_n833_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n830_), .A2(KEYINPUT123), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n820_), .B(new_n839_), .C1(new_n827_), .C2(new_n829_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n638_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n835_), .B1(new_n841_), .B2(new_n792_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n837_), .B1(new_n842_), .B2(new_n833_), .ZN(new_n843_));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n622_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n792_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n836_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT124), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n842_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n622_), .A2(G113gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n844_), .A2(new_n851_), .ZN(G1340gat));
  OAI21_X1  g651(.A(G120gat), .B1(new_n843_), .B2(new_n265_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n265_), .A2(KEYINPUT60), .ZN(new_n854_));
  MUX2_X1   g653(.A(new_n854_), .B(KEYINPUT60), .S(G120gat), .Z(new_n855_));
  NAND3_X1  g654(.A1(new_n847_), .A2(new_n849_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n843_), .B2(new_n638_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n322_), .A2(new_n323_), .A3(G127gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n847_), .A2(new_n849_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1342gat));
  OAI21_X1  g660(.A(G134gat), .B1(new_n843_), .B2(new_n680_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n628_), .A2(G134gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n847_), .A2(new_n849_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1343gat));
  NOR3_X1   g664(.A1(new_n658_), .A2(new_n552_), .A3(new_n499_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n845_), .A2(new_n407_), .A3(new_n699_), .A4(new_n866_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g667(.A1(new_n845_), .A2(new_n407_), .A3(new_n637_), .A4(new_n866_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g669(.A1(new_n845_), .A2(new_n407_), .A3(new_n324_), .A4(new_n866_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  NOR2_X1   g672(.A1(new_n628_), .A2(G162gat), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n845_), .A2(new_n407_), .A3(new_n866_), .A4(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n845_), .A2(new_n407_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n866_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n876_), .A2(new_n680_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(G162gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(G1347gat));
  NOR2_X1   g679(.A1(new_n700_), .A2(new_n553_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n658_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n406_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n792_), .B2(new_n831_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n416_), .B1(new_n885_), .B2(new_n699_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n886_), .A2(KEYINPUT62), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n885_), .A2(new_n448_), .A3(new_n699_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(KEYINPUT62), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(G1348gat));
  AOI21_X1  g689(.A(G176gat), .B1(new_n885_), .B2(new_n637_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n407_), .B1(new_n841_), .B2(new_n792_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n882_), .A2(new_n417_), .A3(new_n265_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(G1349gat));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n883_), .A2(new_n324_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G183gat), .B1(new_n892_), .B2(new_n897_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n319_), .A2(new_n321_), .A3(new_n470_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n885_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n895_), .B1(new_n898_), .B2(new_n901_), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n407_), .B(new_n896_), .C1(new_n841_), .C2(new_n792_), .ZN(new_n903_));
  OAI211_X1 g702(.A(KEYINPUT125), .B(new_n900_), .C1(new_n903_), .C2(G183gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1350gat));
  NAND3_X1  g704(.A1(new_n885_), .A2(new_n629_), .A3(new_n436_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n885_), .A2(new_n679_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n425_), .ZN(G1351gat));
  NAND2_X1  g707(.A1(new_n881_), .A2(new_n560_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n845_), .A2(new_n407_), .A3(new_n699_), .A4(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g711(.A1(new_n845_), .A2(new_n407_), .A3(new_n637_), .A4(new_n910_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g713(.A(new_n638_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n845_), .A2(new_n407_), .A3(new_n910_), .A4(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT126), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n916_), .B(new_n918_), .ZN(G1354gat));
  NOR2_X1   g718(.A1(new_n876_), .A2(new_n909_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n679_), .A2(G218gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n845_), .A2(new_n629_), .A3(new_n407_), .A4(new_n910_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n920_), .A2(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1355gat));
endmodule


