//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT21), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n203_), .B1(KEYINPUT85), .B2(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(KEYINPUT85), .B2(new_n204_), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n207_), .A2(G204gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT84), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT21), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n202_), .B1(new_n210_), .B2(new_n204_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(new_n204_), .B2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n206_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n222_), .B(KEYINPUT83), .Z(new_n223_));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225_));
  OAI22_X1  g024(.A1(new_n224_), .A2(new_n225_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n226_), .B1(new_n225_), .B2(new_n224_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n219_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n224_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n220_), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n218_), .B(KEYINPUT1), .Z(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(new_n217_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n234_));
  OAI21_X1  g033(.A(new_n213_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G228gat), .A3(G233gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G228gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n213_), .B(new_n237_), .C1(new_n233_), .C2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G78gat), .B(G106gat), .Z(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT87), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n241_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n233_), .A2(new_n238_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT28), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G22gat), .B(G50gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n240_), .A2(new_n243_), .A3(new_n241_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n242_), .A2(KEYINPUT88), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n242_), .A2(KEYINPUT88), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(new_n250_), .A4(new_n245_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G127gat), .B(G134gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(G113gat), .B(G120gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n233_), .B(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT4), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n264_), .B(new_n261_), .C1(new_n228_), .C2(new_n232_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT97), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT98), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n262_), .A2(new_n266_), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT99), .Z(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G1gat), .B(G29gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G85gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT0), .B(G57gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n270_), .A2(new_n277_), .A3(new_n272_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n258_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n206_), .A2(new_n212_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284_));
  INV_X1    g083(.A(G169gat), .ZN(new_n285_));
  INV_X1    g084(.A(G176gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT24), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT94), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n284_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(new_n288_), .B2(new_n287_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n291_), .A2(G183gat), .A3(G190gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(G183gat), .B2(G190gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(new_n284_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT26), .B(G190gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(KEYINPUT93), .Z(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT92), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n290_), .B(new_n296_), .C1(new_n298_), .C2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n283_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G169gat), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n293_), .A2(KEYINPUT80), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n293_), .A2(KEYINPUT80), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n292_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n304_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT20), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT102), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n304_), .B1(new_n294_), .B2(new_n308_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n299_), .A2(new_n297_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n284_), .A2(new_n295_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n315_), .B(new_n316_), .C1(new_n284_), .C2(new_n287_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n314_), .B1(new_n307_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n213_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n310_), .A2(KEYINPUT102), .A3(KEYINPUT20), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n313_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT20), .B1(new_n213_), .B2(new_n318_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT91), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n327_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n309_), .B(KEYINPUT95), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n330_), .A2(new_n301_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n328_), .B(new_n329_), .C1(new_n331_), .C2(new_n283_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n324_), .B(KEYINPUT90), .ZN(new_n333_));
  OAI22_X1  g132(.A1(new_n321_), .A2(new_n325_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G8gat), .B(G36gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT18), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n332_), .A2(new_n333_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n302_), .A2(new_n330_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n342_), .A2(KEYINPUT20), .A3(new_n325_), .A4(new_n319_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n338_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(KEYINPUT27), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT103), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n339_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(KEYINPUT96), .A3(new_n350_), .ZN(new_n351_));
  OR3_X1    g150(.A1(new_n345_), .A2(KEYINPUT96), .A3(new_n338_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n340_), .A2(KEYINPUT103), .A3(KEYINPUT27), .A4(new_n346_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n282_), .A2(new_n349_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n263_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n277_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT33), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n280_), .B2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n280_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT101), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT101), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n280_), .A2(new_n366_), .A3(new_n363_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n338_), .A2(KEYINPUT32), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n344_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n334_), .B2(new_n370_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n362_), .A2(new_n368_), .B1(new_n372_), .B2(new_n281_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n356_), .B1(new_n373_), .B2(new_n257_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n261_), .B(KEYINPUT31), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G43gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n318_), .B(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(G15gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT30), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n378_), .B(new_n382_), .Z(new_n383_));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n375_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  OR3_X1    g184(.A1(new_n385_), .A2(new_n384_), .A3(new_n383_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n385_), .B1(new_n384_), .B2(new_n383_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n349_), .A2(new_n354_), .A3(new_n258_), .A4(new_n355_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n281_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n388_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n374_), .A2(new_n388_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G229gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(G1gat), .ZN(new_n397_));
  INV_X1    g196(.A(G8gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT14), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n380_), .A2(KEYINPUT75), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G15gat), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n400_), .A2(new_n402_), .A3(G22gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(G22gat), .B1(new_n400_), .B2(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n399_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G1gat), .B(G8gat), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n406_), .B(new_n399_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G29gat), .B(G36gat), .Z(new_n412_));
  XOR2_X1   g211(.A(G43gat), .B(G50gat), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G29gat), .B(G36gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G43gat), .B(G50gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT77), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(KEYINPUT77), .A3(new_n417_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n411_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n420_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(new_n418_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n410_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n396_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n414_), .A2(KEYINPUT15), .A3(new_n417_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT15), .B1(new_n414_), .B2(new_n417_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n410_), .A3(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT78), .B1(new_n424_), .B2(new_n410_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n429_), .A2(new_n410_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n426_), .B1(new_n434_), .B2(new_n396_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT79), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G113gat), .B(G141gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G169gat), .B(G197gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n442_), .B1(new_n435_), .B2(KEYINPUT79), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G120gat), .B(G148gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT5), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G176gat), .B(G204gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT12), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT70), .ZN(new_n451_));
  INV_X1    g250(.A(G64gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G57gat), .ZN(new_n453_));
  INV_X1    g252(.A(G57gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G64gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT11), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G71gat), .B(G78gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT68), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G71gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G78gat), .ZN(new_n460_));
  INV_X1    g259(.A(G78gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G71gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT68), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G57gat), .B(G64gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n463_), .B(new_n464_), .C1(new_n465_), .C2(KEYINPUT11), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(KEYINPUT11), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n458_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n458_), .B2(new_n466_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n451_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n458_), .A2(new_n466_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n467_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n458_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(KEYINPUT70), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n450_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT6), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n478_), .A2(new_n480_), .A3(KEYINPUT67), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT67), .B1(new_n478_), .B2(new_n480_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT10), .ZN(new_n484_));
  INV_X1    g283(.A(G99gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT64), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n486_), .A2(KEYINPUT64), .A3(new_n487_), .A4(new_n488_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT9), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT66), .B1(G85gat), .B2(G92gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n497_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n494_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT9), .B1(new_n496_), .B2(new_n499_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n483_), .B(new_n493_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n478_), .A2(new_n480_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT67), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n478_), .A2(new_n480_), .A3(KEYINPUT67), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n507_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n497_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n513_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT69), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n478_), .A2(new_n480_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n509_), .A2(new_n510_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n516_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT8), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n520_), .A2(new_n521_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n521_), .B1(new_n520_), .B2(new_n525_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n504_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n476_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n518_), .B1(new_n483_), .B2(new_n511_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n511_), .A2(new_n505_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n517_), .B1(new_n531_), .B2(new_n516_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n504_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n473_), .A2(new_n474_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT12), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G230gat), .A2(G233gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n529_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n536_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n533_), .A2(new_n534_), .ZN(new_n541_));
  OAI211_X1 g340(.A(G230gat), .B(G233gat), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n449_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n539_), .A2(new_n542_), .A3(new_n449_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(KEYINPUT71), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n539_), .A2(new_n542_), .A3(new_n449_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n548_), .B2(new_n543_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT13), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT13), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n395_), .A2(new_n444_), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n528_), .A2(new_n429_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT73), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n528_), .A2(KEYINPUT73), .A3(new_n429_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n533_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n414_), .A2(new_n417_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n564_), .A2(new_n565_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n562_), .A2(new_n563_), .A3(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n562_), .A2(new_n574_), .A3(new_n563_), .A4(new_n570_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n559_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n573_), .A2(KEYINPUT74), .A3(new_n575_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n573_), .A2(KEYINPUT74), .A3(new_n575_), .A4(new_n578_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n576_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AOI211_X1 g383(.A(KEYINPUT37), .B(new_n576_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G127gat), .B(G155gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT16), .ZN(new_n588_));
  XOR2_X1   g387(.A(G183gat), .B(G211gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT76), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n410_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(new_n534_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n471_), .A2(new_n475_), .ZN(new_n600_));
  AOI211_X1 g399(.A(new_n591_), .B(new_n590_), .C1(new_n595_), .C2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n600_), .B2(new_n595_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n586_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n555_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT104), .Z(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n397_), .A3(new_n281_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n608_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n582_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n603_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n555_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n391_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n609_), .A2(new_n610_), .A3(new_n614_), .ZN(G1324gat));
  AND2_X1   g414(.A1(new_n349_), .A2(new_n355_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n354_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G8gat), .B1(new_n613_), .B2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(KEYINPUT105), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT39), .B1(new_n619_), .B2(KEYINPUT105), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n621_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n606_), .A2(new_n398_), .A3(new_n617_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n622_), .A2(KEYINPUT40), .A3(new_n623_), .A4(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  OAI21_X1  g428(.A(G15gat), .B1(new_n613_), .B2(new_n388_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT106), .Z(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT41), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(KEYINPUT41), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n606_), .A2(new_n380_), .A3(new_n392_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(G1326gat));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n606_), .A2(new_n636_), .A3(new_n257_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G22gat), .B1(new_n613_), .B2(new_n258_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1327gat));
  INV_X1    g439(.A(new_n603_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n582_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n555_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n281_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n374_), .A2(new_n388_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n390_), .A2(new_n394_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n586_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(KEYINPUT43), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT108), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n651_));
  INV_X1    g450(.A(new_n649_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n395_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n586_), .B1(new_n395_), .B2(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n645_), .A2(new_n655_), .A3(new_n646_), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT43), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n654_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n554_), .A2(new_n444_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n603_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT44), .B1(new_n659_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  AOI211_X1 g463(.A(new_n664_), .B(new_n661_), .C1(new_n654_), .C2(new_n658_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n281_), .A2(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n644_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n643_), .A2(new_n669_), .A3(new_n617_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT45), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n663_), .A2(new_n665_), .A3(new_n618_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n669_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT46), .B(new_n671_), .C1(new_n672_), .C2(new_n669_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1329gat));
  INV_X1    g476(.A(G43gat), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n388_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n666_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n643_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n681_), .B2(new_n388_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT47), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n680_), .A2(new_n685_), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n643_), .B2(new_n257_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n257_), .A2(G50gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n666_), .B2(new_n689_), .ZN(G1331gat));
  NAND4_X1  g489(.A1(new_n647_), .A2(new_n444_), .A3(new_n554_), .A4(new_n612_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G57gat), .B1(new_n691_), .B2(new_n391_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n647_), .A2(new_n444_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n693_), .A2(KEYINPUT109), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(KEYINPUT109), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(new_n554_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n604_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n281_), .A2(new_n454_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n692_), .B1(new_n697_), .B2(new_n698_), .ZN(G1332gat));
  OAI21_X1  g498(.A(G64gat), .B1(new_n691_), .B2(new_n618_), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n617_), .A2(new_n452_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n697_), .B2(new_n703_), .ZN(G1333gat));
  OAI21_X1  g503(.A(G71gat), .B1(new_n691_), .B2(new_n388_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT49), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n392_), .A2(new_n459_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n697_), .B2(new_n707_), .ZN(G1334gat));
  OAI21_X1  g507(.A(G78gat), .B1(new_n691_), .B2(new_n258_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT50), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n257_), .A2(new_n461_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n697_), .B2(new_n711_), .ZN(G1335gat));
  INV_X1    g511(.A(new_n444_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n641_), .A2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n659_), .A2(new_n554_), .A3(new_n281_), .A4(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(G85gat), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n694_), .A2(new_n554_), .A3(new_n642_), .A4(new_n695_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n717_), .A2(G85gat), .A3(new_n391_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1336gat));
  INV_X1    g520(.A(new_n659_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n554_), .A2(new_n714_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n722_), .A2(new_n618_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(G92gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n617_), .A2(new_n725_), .ZN(new_n726_));
  OAI22_X1  g525(.A1(new_n724_), .A2(new_n725_), .B1(new_n717_), .B2(new_n726_), .ZN(G1337gat));
  NOR2_X1   g526(.A1(new_n722_), .A2(new_n723_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n485_), .B1(new_n728_), .B2(new_n392_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n392_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT112), .B1(new_n717_), .B2(new_n730_), .ZN(new_n731_));
  OR3_X1    g530(.A1(new_n729_), .A2(KEYINPUT51), .A3(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT51), .B1(new_n729_), .B2(new_n731_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1338gat));
  NAND4_X1  g533(.A1(new_n659_), .A2(new_n554_), .A3(new_n257_), .A4(new_n714_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G106gat), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n258_), .A2(G106gat), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n696_), .A2(new_n739_), .A3(new_n642_), .A4(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n740_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT113), .B1(new_n717_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n735_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n738_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n738_), .A2(new_n744_), .A3(new_n748_), .A4(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  NOR2_X1   g549(.A1(new_n554_), .A2(new_n713_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n604_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT54), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n604_), .A2(new_n751_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n538_), .B1(new_n529_), .B2(new_n537_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n539_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n529_), .A2(new_n537_), .A3(KEYINPUT55), .A4(new_n538_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n761_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n448_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n441_), .A2(new_n443_), .A3(new_n545_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT56), .B1(new_n761_), .B2(new_n448_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n766_), .B(new_n449_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n396_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n431_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n422_), .A2(new_n425_), .A3(new_n396_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n440_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n546_), .A2(new_n549_), .A3(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT57), .B(new_n582_), .C1(new_n770_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778_));
  INV_X1    g577(.A(new_n426_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n429_), .A2(new_n410_), .A3(new_n430_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n430_), .B1(new_n411_), .B2(new_n421_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n429_), .A2(new_n410_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n779_), .B(new_n440_), .C1(new_n783_), .C2(new_n771_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n772_), .A2(new_n773_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n440_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n778_), .B1(new_n786_), .B2(new_n548_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n775_), .A2(KEYINPUT116), .A3(new_n545_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI221_X1 g591(.A(new_n789_), .B1(KEYINPUT117), .B2(KEYINPUT58), .C1(new_n765_), .C2(new_n767_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n792_), .B(new_n793_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n777_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n582_), .B1(new_n770_), .B2(new_n776_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n795_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n756_), .B1(new_n641_), .B2(new_n798_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n389_), .A2(new_n388_), .A3(new_n391_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n799_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n761_), .A2(new_n448_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n766_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n448_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n769_), .A3(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n762_), .A2(new_n763_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n776_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n796_), .B1(new_n808_), .B2(new_n611_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT115), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n797_), .A2(new_n811_), .A3(new_n796_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n795_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n603_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n777_), .A2(new_n794_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n811_), .B1(new_n797_), .B2(new_n796_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n776_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n765_), .A2(new_n767_), .A3(KEYINPUT114), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n764_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT115), .B(KEYINPUT57), .C1(new_n820_), .C2(new_n582_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n816_), .B(new_n814_), .C1(new_n817_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n756_), .B(KEYINPUT119), .C1(new_n815_), .C2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n816_), .B1(new_n817_), .B2(new_n821_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT118), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n603_), .A3(new_n822_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT119), .B1(new_n828_), .B2(new_n756_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n825_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n800_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n802_), .B1(new_n831_), .B2(KEYINPUT59), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n832_), .A2(new_n713_), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n713_), .A2(new_n834_), .ZN(new_n835_));
  OAI22_X1  g634(.A1(new_n833_), .A2(new_n834_), .B1(new_n831_), .B2(new_n835_), .ZN(G1340gat));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n837_));
  AOI21_X1  g636(.A(G120gat), .B1(new_n554_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT60), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n831_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n832_), .A2(new_n554_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n839_), .B2(new_n844_), .ZN(G1341gat));
  AND2_X1   g644(.A1(new_n832_), .A2(new_n641_), .ZN(new_n846_));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n641_), .A2(new_n847_), .ZN(new_n848_));
  OAI22_X1  g647(.A1(new_n846_), .A2(new_n847_), .B1(new_n831_), .B2(new_n848_), .ZN(G1342gat));
  AND2_X1   g648(.A1(new_n832_), .A2(new_n586_), .ZN(new_n850_));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n611_), .A2(new_n851_), .ZN(new_n852_));
  OAI22_X1  g651(.A1(new_n850_), .A2(new_n851_), .B1(new_n831_), .B2(new_n852_), .ZN(G1343gat));
  NOR3_X1   g652(.A1(new_n617_), .A2(new_n391_), .A3(new_n258_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n830_), .A2(KEYINPUT121), .A3(new_n388_), .A4(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n756_), .B1(new_n815_), .B2(new_n823_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n858_), .A2(new_n388_), .A3(new_n824_), .A4(new_n854_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n855_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n713_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n554_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n862_), .B2(new_n641_), .ZN(new_n868_));
  AOI211_X1 g667(.A(KEYINPUT122), .B(new_n603_), .C1(new_n855_), .C2(new_n861_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n868_), .A2(new_n869_), .A3(new_n871_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n859_), .A2(new_n860_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n859_), .A2(new_n860_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n641_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT122), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n862_), .A2(new_n867_), .A3(new_n641_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n870_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n872_), .A2(new_n878_), .ZN(G1346gat));
  INV_X1    g678(.A(new_n862_), .ZN(new_n880_));
  OR3_X1    g679(.A1(new_n880_), .A2(G162gat), .A3(new_n582_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G162gat), .B1(new_n880_), .B2(new_n648_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1347gat));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n618_), .A2(new_n393_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n799_), .A2(new_n258_), .A3(new_n885_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n886_), .A2(new_n713_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT22), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n884_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G169gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n285_), .B1(new_n887_), .B2(new_n884_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n889_), .B2(new_n891_), .ZN(G1348gat));
  AOI21_X1  g691(.A(G176gat), .B1(new_n886_), .B2(new_n554_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n830_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n257_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n885_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n896_), .A2(new_n286_), .A3(new_n553_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n893_), .B1(new_n895_), .B2(new_n897_), .ZN(G1349gat));
  NAND3_X1  g697(.A1(new_n886_), .A2(new_n300_), .A3(new_n641_), .ZN(new_n899_));
  NOR4_X1   g698(.A1(new_n894_), .A2(new_n257_), .A3(new_n603_), .A4(new_n896_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(G183gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT123), .ZN(G1350gat));
  INV_X1    g701(.A(G190gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n886_), .B2(new_n586_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT124), .ZN(new_n905_));
  INV_X1    g704(.A(new_n298_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n886_), .A2(new_n906_), .A3(new_n611_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1351gat));
  NAND4_X1  g707(.A1(new_n830_), .A2(new_n388_), .A3(new_n282_), .A4(new_n617_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n444_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n207_), .ZN(G1352gat));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n553_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT125), .B(G204gat), .Z(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n912_), .B2(new_n915_), .ZN(G1353gat));
  OR2_X1    g715(.A1(new_n909_), .A2(new_n603_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT63), .B(G211gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n920_));
  INV_X1    g719(.A(G211gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n917_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n917_), .A2(KEYINPUT126), .A3(new_n920_), .A4(new_n921_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n919_), .B1(new_n924_), .B2(new_n925_), .ZN(G1354gat));
  INV_X1    g725(.A(G218gat), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n909_), .A2(new_n927_), .A3(new_n648_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n909_), .A2(KEYINPUT127), .A3(new_n582_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(G218gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(KEYINPUT127), .B1(new_n909_), .B2(new_n582_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n928_), .B1(new_n930_), .B2(new_n931_), .ZN(G1355gat));
endmodule


