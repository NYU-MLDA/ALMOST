//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202_));
  OR2_X1    g001(.A1(G197gat), .A2(G204gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT21), .A3(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206_));
  OR3_X1    g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT88), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT88), .B1(new_n205_), .B2(new_n206_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n203_), .A2(new_n204_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT21), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n205_), .A2(new_n206_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G228gat), .A2(G233gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT82), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(KEYINPUT82), .B(new_n224_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n234_));
  OAI22_X1  g033(.A1(new_n224_), .A2(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT83), .ZN(new_n236_));
  INV_X1    g035(.A(new_n233_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n236_), .B1(new_n237_), .B2(KEYINPUT2), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(KEYINPUT83), .A3(new_n234_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n235_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n231_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n231_), .A2(new_n240_), .A3(KEYINPUT84), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n223_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n221_), .B1(KEYINPUT1), .B2(new_n219_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n219_), .A2(KEYINPUT1), .ZN(new_n247_));
  AOI211_X1 g046(.A(new_n224_), .B(new_n237_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n218_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n244_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT84), .B1(new_n231_), .B2(new_n240_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n222_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n248_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT85), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT29), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT87), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n249_), .A2(new_n254_), .A3(new_n258_), .A4(KEYINPUT29), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n217_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n215_), .B1(new_n262_), .B2(new_n214_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G78gat), .B(G106gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n202_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G22gat), .B(G50gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT28), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT86), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n255_), .A2(new_n271_), .A3(new_n256_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n271_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n270_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n272_), .A3(new_n269_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n265_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n260_), .A2(new_n265_), .A3(new_n263_), .ZN(new_n281_));
  OAI22_X1  g080(.A1(new_n267_), .A2(new_n278_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n278_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n202_), .A4(new_n279_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT20), .ZN(new_n287_));
  NOR3_X1   g086(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT25), .B(G183gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT24), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(G169gat), .B2(G176gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(G169gat), .B2(G176gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(G183gat), .B2(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT78), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(G183gat), .A3(G190gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n297_), .B1(new_n302_), .B2(new_n296_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n295_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n296_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT79), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G169gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n304_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n287_), .B1(new_n314_), .B2(new_n214_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT19), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n305_), .A2(new_n307_), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n293_), .A2(KEYINPUT91), .B1(G169gat), .B2(G176gat), .ZN(new_n320_));
  INV_X1    g119(.A(G169gat), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT24), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT91), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n319_), .B(new_n291_), .C1(new_n320_), .C2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n312_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n315_), .B(new_n318_), .C1(new_n214_), .C2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT18), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  AOI21_X1  g132(.A(new_n287_), .B1(new_n328_), .B2(new_n214_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n207_), .A2(new_n208_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n335_), .B(new_n304_), .C1(new_n310_), .C2(new_n313_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n318_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT92), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AOI211_X1 g138(.A(KEYINPUT92), .B(new_n318_), .C1(new_n334_), .C2(new_n336_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n329_), .B(new_n333_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n333_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n214_), .B1(new_n328_), .B2(KEYINPUT97), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(KEYINPUT97), .B2(new_n328_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n318_), .B1(new_n344_), .B2(new_n315_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n334_), .A2(new_n336_), .A3(new_n318_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n342_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n341_), .A2(new_n347_), .A3(KEYINPUT27), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n337_), .B(new_n338_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(KEYINPUT93), .A3(new_n333_), .A4(new_n329_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT93), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n341_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n329_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n342_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n348_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n286_), .A2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G1gat), .B(G29gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G113gat), .B(G120gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND3_X1  g168(.A1(new_n249_), .A2(new_n254_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OR3_X1    g172(.A1(new_n245_), .A2(new_n248_), .A3(new_n369_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n366_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT95), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n370_), .A2(new_n374_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n366_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n370_), .A2(new_n374_), .A3(KEYINPUT95), .A4(new_n365_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n364_), .B1(new_n377_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n364_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n376_), .A2(new_n384_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(G71gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G99gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n314_), .B(new_n391_), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(new_n369_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G15gat), .B(G43gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT80), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT30), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT31), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n393_), .B(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n386_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n359_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n386_), .ZN(new_n401_));
  AND4_X1   g200(.A1(new_n401_), .A2(new_n282_), .A3(new_n285_), .A4(new_n357_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n364_), .B1(new_n379_), .B2(new_n365_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n375_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n372_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n405_), .B2(new_n365_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(new_n355_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n385_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n382_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n410_), .A2(KEYINPUT33), .A3(new_n384_), .A4(new_n376_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT96), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n407_), .A2(new_n409_), .A3(new_n411_), .A4(KEYINPUT96), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n345_), .A2(new_n346_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n333_), .A2(KEYINPUT32), .ZN(new_n417_));
  MUX2_X1   g216(.A(new_n416_), .B(new_n353_), .S(new_n417_), .Z(new_n418_));
  NAND2_X1  g217(.A1(new_n386_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(new_n415_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n286_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n402_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n398_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n400_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G232gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT34), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT35), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n430_), .A2(KEYINPUT70), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT65), .ZN(new_n432_));
  INV_X1    g231(.A(G106gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n390_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT7), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G99gat), .A2(G106gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT6), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(G99gat), .A3(G106gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT7), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n432_), .A2(new_n441_), .A3(new_n390_), .A4(new_n433_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n435_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(G85gat), .ZN(new_n444_));
  INV_X1    g243(.A(G92gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G85gat), .A2(G92gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT8), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n443_), .A2(new_n453_), .A3(new_n449_), .ZN(new_n456_));
  OR2_X1    g255(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n433_), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n446_), .A2(KEYINPUT9), .A3(new_n447_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n447_), .A2(KEYINPUT9), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n440_), .A2(new_n459_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n455_), .A2(new_n456_), .A3(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G29gat), .B(G36gat), .Z(new_n464_));
  XOR2_X1   g263(.A(G43gat), .B(G50gat), .Z(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n463_), .A2(new_n466_), .B1(new_n428_), .B2(new_n427_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT69), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n464_), .B(new_n465_), .Z(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT15), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  AND4_X1   g272(.A1(new_n440_), .A2(new_n459_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(new_n454_), .B2(new_n450_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n456_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n468_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  AND4_X1   g276(.A1(new_n468_), .A2(new_n476_), .A3(new_n470_), .A4(new_n472_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n467_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n430_), .A2(KEYINPUT70), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n431_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(new_n431_), .A3(new_n480_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G190gat), .B(G218gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G134gat), .B(G162gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT36), .Z(new_n487_));
  NAND3_X1  g286(.A1(new_n482_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n486_), .A2(KEYINPUT36), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n479_), .A2(new_n431_), .A3(new_n480_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(new_n490_), .B2(new_n481_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT71), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n488_), .A2(new_n491_), .A3(new_n492_), .A4(KEYINPUT37), .ZN(new_n496_));
  XOR2_X1   g295(.A(G127gat), .B(G155gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT16), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G183gat), .B(G211gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT72), .B(G1gat), .ZN(new_n501_));
  INV_X1    g300(.A(G8gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT14), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G8gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n512_));
  XOR2_X1   g311(.A(G71gat), .B(G78gat), .Z(new_n513_));
  OR2_X1    g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n513_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n510_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT73), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n518_), .B(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n500_), .B1(new_n521_), .B2(KEYINPUT74), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT17), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n521_), .B2(new_n500_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n495_), .A2(new_n496_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n515_), .A2(new_n516_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n512_), .A2(new_n513_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n476_), .A2(new_n531_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n437_), .A2(new_n439_), .B1(new_n533_), .B2(new_n441_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n448_), .B1(new_n534_), .B2(new_n435_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n462_), .B1(new_n535_), .B2(new_n453_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n456_), .ZN(new_n537_));
  OAI211_X1 g336(.A(KEYINPUT12), .B(new_n531_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n476_), .A2(KEYINPUT67), .A3(KEYINPUT12), .A4(new_n531_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n532_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n517_), .B1(new_n475_), .B2(new_n456_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(KEYINPUT12), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT12), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT68), .B(new_n546_), .C1(new_n463_), .C2(new_n517_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT64), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n532_), .B2(new_n544_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G120gat), .B(G148gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G176gat), .B(G204gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n552_), .A2(new_n553_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(KEYINPUT13), .A3(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n528_), .A2(KEYINPUT75), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT75), .B1(new_n528_), .B2(new_n567_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT77), .ZN(new_n570_));
  INV_X1    g369(.A(new_n510_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n510_), .A2(new_n466_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT76), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n572_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n469_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n577_), .B2(new_n573_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G169gat), .B(G197gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n576_), .A2(new_n578_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n577_), .A2(new_n573_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n574_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n572_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n581_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n570_), .B1(new_n583_), .B2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n582_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n587_), .A3(new_n581_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(KEYINPUT77), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n568_), .A2(new_n569_), .A3(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n424_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n386_), .A3(new_n501_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT38), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT98), .Z(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n598_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT99), .Z(new_n602_));
  NOR2_X1   g401(.A1(new_n566_), .A2(new_n594_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n488_), .A2(new_n491_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n526_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n424_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n401_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n602_), .A3(new_n609_), .ZN(G1324gat));
  NAND3_X1  g409(.A1(new_n607_), .A2(KEYINPUT101), .A3(new_n358_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n611_), .A2(G8gat), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n358_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n615_), .A2(new_n611_), .A3(KEYINPUT39), .A4(G8gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n596_), .A2(new_n502_), .A3(new_n358_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n618_), .A2(KEYINPUT40), .A3(new_n619_), .A4(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n619_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT39), .B1(new_n612_), .B2(new_n615_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n623_), .A2(new_n627_), .ZN(G1325gat));
  INV_X1    g427(.A(G15gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n607_), .B2(new_n423_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n596_), .A2(new_n629_), .A3(new_n423_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n286_), .B(KEYINPUT102), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n607_), .B2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT42), .Z(new_n638_));
  NAND3_X1  g437(.A1(new_n596_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1327gat));
  INV_X1    g439(.A(new_n603_), .ZN(new_n641_));
  AOI22_X1  g440(.A1(new_n412_), .A2(new_n413_), .B1(new_n386_), .B2(new_n418_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n286_), .B1(new_n642_), .B2(new_n415_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n398_), .B1(new_n643_), .B2(new_n402_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n641_), .B1(new_n644_), .B2(new_n400_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n604_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n526_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n648_), .A2(G29gat), .A3(new_n401_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n641_), .A2(new_n526_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n495_), .A2(new_n496_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT43), .B(new_n652_), .C1(new_n644_), .C2(new_n400_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n424_), .B2(new_n651_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n650_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(KEYINPUT44), .B(new_n650_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n386_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(G29gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n660_), .B2(G29gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n649_), .B1(new_n662_), .B2(new_n663_), .ZN(G1328gat));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n658_), .A2(new_n358_), .A3(new_n659_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G36gat), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n357_), .A2(G36gat), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n424_), .A2(new_n603_), .A3(new_n647_), .A4(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n645_), .A2(new_n647_), .A3(new_n673_), .A4(new_n671_), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n675_), .A2(new_n676_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n668_), .B1(new_n670_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n677_), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n667_), .B(new_n679_), .C1(new_n669_), .C2(G36gat), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1329gat));
  NAND4_X1  g480(.A1(new_n658_), .A2(G43gat), .A3(new_n423_), .A4(new_n659_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n424_), .A2(new_n423_), .A3(new_n603_), .A4(new_n647_), .ZN(new_n683_));
  INV_X1    g482(.A(G43gat), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT106), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n682_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g487(.A1(new_n658_), .A2(G50gat), .A3(new_n286_), .A4(new_n659_), .ZN(new_n689_));
  INV_X1    g488(.A(G50gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(new_n648_), .B2(new_n635_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1331gat));
  AOI211_X1 g491(.A(new_n567_), .B(new_n593_), .C1(new_n644_), .C2(new_n400_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(new_n606_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n401_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n693_), .A2(new_n528_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n386_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1332gat));
  NOR2_X1   g499(.A1(new_n357_), .A2(G64gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT107), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n697_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G64gat), .B1(new_n695_), .B2(new_n357_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT48), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT48), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(G1333gat));
  AOI21_X1  g506(.A(new_n388_), .B1(new_n694_), .B2(new_n423_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT49), .Z(new_n709_));
  NOR2_X1   g508(.A1(new_n398_), .A2(G71gat), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT108), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n697_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1334gat));
  INV_X1    g512(.A(G78gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n694_), .B2(new_n636_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT50), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n697_), .A2(new_n714_), .A3(new_n636_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1335gat));
  OR2_X1    g517(.A1(new_n653_), .A2(new_n655_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n567_), .A2(new_n526_), .A3(new_n593_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n444_), .B1(new_n721_), .B2(new_n386_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n693_), .A2(new_n647_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n723_), .A2(new_n444_), .A3(new_n386_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1336gat));
  NAND3_X1  g524(.A1(new_n723_), .A2(new_n445_), .A3(new_n358_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n721_), .A2(new_n358_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n726_), .B1(new_n728_), .B2(new_n445_), .ZN(G1337gat));
  AND3_X1   g528(.A1(new_n423_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT110), .B1(new_n723_), .B2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n423_), .B(new_n720_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(G99gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G99gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT51), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n738_), .B(new_n731_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1338gat));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n286_), .B(new_n720_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n743_), .B2(new_n433_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n693_), .A2(new_n433_), .A3(new_n286_), .A4(new_n647_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT111), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT53), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n744_), .A2(new_n746_), .A3(new_n750_), .A4(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1339gat));
  NAND3_X1  g551(.A1(new_n528_), .A2(new_n567_), .A3(new_n594_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(KEYINPUT112), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n753_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT118), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n593_), .A2(new_n561_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n551_), .B1(new_n542_), .B2(new_n548_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n552_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n542_), .A2(new_n548_), .A3(KEYINPUT55), .A4(new_n551_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT56), .B1(new_n766_), .B2(new_n558_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n768_), .B(new_n560_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n761_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT113), .B(new_n761_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n572_), .A2(new_n573_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n575_), .B1(new_n774_), .B2(KEYINPUT114), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(KEYINPUT114), .B2(new_n774_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n581_), .B1(new_n584_), .B2(new_n575_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n583_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n562_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n772_), .A2(new_n773_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n604_), .A2(new_n782_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n780_), .A2(new_n781_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n781_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n778_), .A2(new_n561_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(KEYINPUT115), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(KEYINPUT115), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n787_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n651_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n780_), .A2(new_n646_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n782_), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n760_), .B(new_n526_), .C1(new_n786_), .C2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n782_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n780_), .A2(new_n783_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT116), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n780_), .A2(new_n781_), .A3(new_n783_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n798_), .A2(new_n800_), .A3(new_n793_), .A4(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT118), .B1(new_n802_), .B2(new_n605_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n759_), .B1(new_n797_), .B2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n401_), .A2(new_n398_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n359_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n807_));
  INV_X1    g606(.A(new_n806_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n526_), .B1(new_n786_), .B2(new_n796_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n758_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n804_), .A2(new_n807_), .B1(KEYINPUT59), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n594_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(KEYINPUT117), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n770_), .A2(new_n771_), .B1(new_n562_), .B2(new_n778_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n604_), .B1(new_n815_), .B2(new_n773_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n793_), .B1(new_n816_), .B2(KEYINPUT57), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n817_), .A2(new_n785_), .A3(new_n784_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n759_), .B1(new_n818_), .B2(new_n526_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n808_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n814_), .A2(new_n821_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n594_), .A2(G113gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n813_), .B1(new_n822_), .B2(new_n823_), .ZN(G1340gat));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n811_), .B2(new_n566_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT60), .ZN(new_n828_));
  AOI21_X1  g627(.A(G120gat), .B1(new_n566_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n828_), .B2(G120gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n814_), .A2(new_n821_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n825_), .B1(new_n827_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n810_), .A2(KEYINPUT59), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n760_), .B1(new_n818_), .B2(new_n526_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n802_), .A2(KEYINPUT118), .A3(new_n605_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n758_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n807_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n566_), .B(new_n834_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(G120gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(KEYINPUT119), .A3(new_n831_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n833_), .A2(new_n841_), .ZN(G1341gat));
  NAND3_X1  g641(.A1(new_n814_), .A2(new_n526_), .A3(new_n821_), .ZN(new_n843_));
  INV_X1    g642(.A(G127gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(KEYINPUT120), .A3(new_n844_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n605_), .A2(new_n844_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n847_), .A2(new_n848_), .B1(new_n811_), .B2(new_n849_), .ZN(G1342gat));
  NAND3_X1  g649(.A1(new_n814_), .A2(new_n604_), .A3(new_n821_), .ZN(new_n851_));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n651_), .A2(G134gat), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT121), .Z(new_n855_));
  OAI211_X1 g654(.A(new_n834_), .B(new_n855_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n853_), .A2(KEYINPUT122), .A3(new_n856_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1343gat));
  NOR4_X1   g660(.A1(new_n421_), .A2(new_n358_), .A3(new_n401_), .A4(new_n423_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n819_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n594_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT123), .B(G141gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n863_), .A2(new_n567_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g667(.A1(new_n863_), .A2(new_n605_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT61), .B(G155gat), .Z(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n863_), .B2(new_n652_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n646_), .A2(G162gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n863_), .B2(new_n873_), .ZN(G1347gat));
  NAND2_X1  g673(.A1(new_n399_), .A2(new_n358_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n635_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n837_), .A2(new_n877_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT22), .B(G169gat), .Z(new_n879_));
  NOR2_X1   g678(.A1(new_n594_), .A2(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT125), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  INV_X1    g682(.A(new_n877_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n593_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n835_), .A2(new_n836_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n759_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n321_), .B1(new_n887_), .B2(KEYINPUT124), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n837_), .B2(new_n885_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n883_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n804_), .A2(KEYINPUT124), .A3(new_n593_), .A4(new_n884_), .ZN(new_n892_));
  AND4_X1   g691(.A1(new_n883_), .A2(new_n890_), .A3(new_n892_), .A4(G169gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n882_), .B1(new_n891_), .B2(new_n893_), .ZN(G1348gat));
  AOI21_X1  g693(.A(G176gat), .B1(new_n878_), .B2(new_n566_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n758_), .B1(new_n802_), .B2(new_n605_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n286_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n875_), .A2(new_n322_), .A3(new_n567_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n897_), .B2(new_n898_), .ZN(G1349gat));
  NOR2_X1   g698(.A1(new_n875_), .A2(new_n605_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G183gat), .B1(new_n897_), .B2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n605_), .A2(new_n289_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n878_), .B2(new_n902_), .ZN(G1350gat));
  INV_X1    g702(.A(new_n878_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G190gat), .B1(new_n904_), .B2(new_n652_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n878_), .A2(new_n290_), .A3(new_n604_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1351gat));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n286_), .A2(new_n401_), .A3(new_n358_), .A4(new_n398_), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n896_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n896_), .B2(new_n909_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n593_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n566_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AND4_X1   g717(.A1(new_n526_), .A2(new_n912_), .A3(new_n917_), .A4(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n912_), .B2(new_n526_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1354gat));
  INV_X1    g720(.A(G218gat), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n912_), .B2(new_n651_), .ZN(new_n923_));
  AOI211_X1 g722(.A(G218gat), .B(new_n646_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT127), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n912_), .A2(new_n922_), .A3(new_n604_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n652_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n926_), .B(new_n927_), .C1(new_n922_), .C2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n929_), .ZN(G1355gat));
endmodule


