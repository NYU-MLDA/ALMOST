//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT86), .ZN(new_n203_));
  XOR2_X1   g002(.A(G15gat), .B(G43gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT82), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT82), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G169gat), .A3(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT22), .B(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n216_), .B(new_n217_), .C1(G183gat), .C2(G190gat), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n210_), .A2(new_n213_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT26), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT80), .B1(new_n222_), .B2(G190gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n229_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT80), .B1(new_n221_), .B2(new_n223_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT81), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n212_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n210_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n219_), .B1(new_n234_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT30), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(KEYINPUT30), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n204_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n204_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n243_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT83), .B(KEYINPUT84), .Z(new_n251_));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G71gat), .B(G99gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n253_), .B(new_n254_), .Z(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n250_), .A2(new_n256_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n203_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n259_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(KEYINPUT86), .A3(new_n257_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G127gat), .B(G134gat), .Z(new_n263_));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G127gat), .B(G134gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT85), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G113gat), .B(G120gat), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n265_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n268_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT31), .Z(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(new_n262_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n272_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n203_), .B(new_n274_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT97), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT19), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G204gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n282_), .B1(KEYINPUT91), .B2(G197gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT90), .B(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(G197gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(KEYINPUT91), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n283_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT21), .ZN(new_n288_));
  NOR2_X1   g087(.A1(KEYINPUT91), .A2(KEYINPUT21), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(KEYINPUT90), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G204gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n285_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n289_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n288_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n298_), .A2(KEYINPUT21), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n293_), .A2(new_n294_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n238_), .B1(new_n205_), .B2(new_n240_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT92), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n224_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n221_), .A2(new_n223_), .A3(KEYINPUT92), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(new_n228_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n209_), .B1(new_n212_), .B2(new_n211_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n218_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT20), .B1(new_n302_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n234_), .A2(new_n241_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n310_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT95), .B1(new_n315_), .B2(new_n302_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n298_), .B1(new_n287_), .B2(KEYINPUT21), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n317_), .A2(new_n295_), .B1(new_n300_), .B2(new_n299_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT95), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n242_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n281_), .B(new_n313_), .C1(new_n316_), .C2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT96), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n315_), .A2(KEYINPUT95), .A3(new_n302_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n319_), .B1(new_n242_), .B2(new_n318_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n312_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT96), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n281_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(new_n242_), .B2(new_n318_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n303_), .A2(new_n307_), .B1(new_n309_), .B2(new_n218_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n318_), .A2(new_n330_), .A3(KEYINPUT93), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT93), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n302_), .B2(new_n311_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n329_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n334_), .A2(KEYINPUT94), .A3(new_n280_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT94), .B1(new_n334_), .B2(new_n280_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n322_), .B(new_n327_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT18), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n278_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n322_), .A2(new_n327_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n334_), .A2(new_n280_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n334_), .A2(KEYINPUT94), .A3(new_n280_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n344_), .A2(KEYINPUT97), .A3(new_n349_), .A4(new_n341_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n337_), .A2(new_n342_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n343_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  INV_X1    g154(.A(G141gat), .ZN(new_n356_));
  INV_X1    g155(.A(G148gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT1), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT88), .ZN(new_n361_));
  OR3_X1    g160(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n362_), .B(new_n363_), .C1(KEYINPUT1), .C2(new_n359_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n355_), .B(new_n358_), .C1(new_n361_), .C2(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n362_), .A2(new_n363_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n358_), .A2(KEYINPUT3), .ZN(new_n367_));
  OR3_X1    g166(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT89), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n369_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(KEYINPUT2), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n367_), .B(new_n368_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n370_), .A2(new_n371_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n359_), .B(new_n366_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n365_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(KEYINPUT29), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n375_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n318_), .B1(KEYINPUT29), .B2(new_n375_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G78gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G106gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G22gat), .B(G50gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n382_), .B(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n375_), .A2(new_n271_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n365_), .B(new_n374_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(KEYINPUT4), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n375_), .A2(new_n271_), .A3(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n389_), .A2(new_n392_), .A3(new_n390_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT98), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G85gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT0), .B(G57gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  NAND4_X1  g202(.A1(new_n389_), .A2(KEYINPUT98), .A3(new_n390_), .A4(new_n392_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n396_), .A2(new_n399_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(KEYINPUT100), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(KEYINPUT100), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n396_), .A2(new_n399_), .A3(new_n404_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n403_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n388_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n337_), .A2(new_n342_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n329_), .B(new_n281_), .C1(new_n331_), .C2(new_n333_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(new_n325_), .B2(new_n281_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT27), .B1(new_n416_), .B2(new_n341_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n354_), .A2(new_n412_), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n389_), .A2(new_n393_), .A3(new_n390_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n409_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n391_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT99), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT99), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n391_), .A2(new_n425_), .A3(new_n392_), .A4(new_n395_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n422_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n399_), .A2(new_n404_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n403_), .A4(new_n396_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n405_), .A2(KEYINPUT33), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n343_), .A2(new_n350_), .A3(new_n351_), .A4(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n415_), .A2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n411_), .B(new_n435_), .C1(new_n337_), .C2(new_n434_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n388_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n277_), .B1(new_n420_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n411_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n273_), .A2(new_n440_), .A3(new_n275_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n418_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(new_n388_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G85gat), .B(G92gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n446_), .A2(KEYINPUT9), .ZN(new_n447_));
  INV_X1    g246(.A(G92gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(KEYINPUT9), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT64), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G99gat), .A2(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT6), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(G99gat), .A3(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT64), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n447_), .A2(new_n449_), .A3(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT10), .B(G99gat), .Z(new_n459_));
  INV_X1    g258(.A(G106gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n451_), .A2(new_n456_), .A3(new_n458_), .A4(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT67), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n453_), .A2(new_n455_), .A3(KEYINPUT66), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT66), .B1(new_n453_), .B2(new_n455_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT66), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n454_), .B1(G99gat), .B2(G106gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n452_), .A2(KEYINPUT6), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n453_), .A2(new_n455_), .A3(KEYINPUT66), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT67), .A3(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT7), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n467_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n446_), .B(KEYINPUT65), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n463_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n456_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n477_), .A2(new_n463_), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n462_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G29gat), .B(G36gat), .Z(new_n482_));
  XOR2_X1   g281(.A(G43gat), .B(G50gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT15), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G232gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT34), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n488_), .A2(KEYINPUT35), .ZN(new_n489_));
  INV_X1    g288(.A(new_n484_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n486_), .B(new_n489_), .C1(new_n490_), .C2(new_n481_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(KEYINPUT35), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT70), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n491_), .B(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G190gat), .B(G218gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT71), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G134gat), .B(G162gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT36), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(KEYINPUT36), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n494_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT101), .Z(new_n504_));
  XNOR2_X1  g303(.A(G57gat), .B(G64gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT11), .ZN(new_n506_));
  XOR2_X1   g305(.A(G71gat), .B(G78gat), .Z(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n505_), .A2(KEYINPUT11), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n506_), .A2(new_n507_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G231gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G8gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n516_), .A2(KEYINPUT73), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(KEYINPUT73), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G1gat), .B(G8gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT74), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n522_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n514_), .B(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n529_));
  NOR2_X1   g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G127gat), .B(G155gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT16), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G183gat), .B(G211gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n528_), .B1(new_n530_), .B2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n534_), .B2(new_n530_), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT77), .Z(new_n537_));
  NOR3_X1   g336(.A1(new_n445_), .A2(new_n504_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n525_), .B(new_n484_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT78), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n485_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n525_), .A2(new_n484_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n540_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT79), .Z(new_n547_));
  NOR2_X1   g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G169gat), .B(G197gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n548_), .B(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n462_), .B(new_n512_), .C1(new_n478_), .C2(new_n480_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(KEYINPUT68), .A3(new_n554_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT12), .ZN(new_n559_));
  INV_X1    g358(.A(new_n512_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n481_), .B2(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n481_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n557_), .B(new_n558_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n481_), .A2(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n553_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(G230gat), .A3(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT5), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G176gat), .B(G204gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n563_), .A2(new_n566_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT69), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n571_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(new_n574_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT13), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n538_), .A2(new_n552_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT102), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n202_), .B1(new_n584_), .B2(new_n411_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n552_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n445_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n503_), .B2(KEYINPUT72), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT72), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n500_), .A2(new_n590_), .A3(KEYINPUT37), .A4(new_n502_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n537_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n582_), .A3(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n594_), .A2(G1gat), .A3(new_n440_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT38), .ZN(new_n596_));
  OR3_X1    g395(.A1(new_n585_), .A2(new_n596_), .A3(KEYINPUT103), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT103), .B1(new_n585_), .B2(new_n596_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(G1324gat));
  OAI21_X1  g398(.A(G8gat), .B1(new_n583_), .B2(new_n442_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT39), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n594_), .A2(G8gat), .A3(new_n442_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT104), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n601_), .A2(KEYINPUT40), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1325gat));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n583_), .B(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G15gat), .B1(new_n611_), .B2(new_n276_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n594_), .A2(G15gat), .A3(new_n276_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT105), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(G1326gat));
  OR3_X1    g416(.A1(new_n594_), .A2(G22gat), .A3(new_n388_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n388_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n584_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT42), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n620_), .A2(new_n621_), .A3(G22gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n620_), .B2(G22gat), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n622_), .B2(new_n623_), .ZN(G1327gat));
  OAI21_X1  g423(.A(new_n592_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT43), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT43), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n627_), .B(new_n592_), .C1(new_n439_), .C2(new_n444_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n582_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n536_), .B(KEYINPUT77), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n630_), .A2(new_n586_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT44), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n629_), .A2(KEYINPUT44), .A3(new_n632_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n411_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G29gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n504_), .A2(new_n537_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n630_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n587_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n440_), .A2(G29gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT106), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n639_), .B1(new_n642_), .B2(new_n644_), .ZN(G1328gat));
  INV_X1    g444(.A(new_n642_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n442_), .A2(G36gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(KEYINPUT45), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT45), .ZN(new_n649_));
  INV_X1    g448(.A(new_n647_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n642_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n442_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n635_), .A2(new_n653_), .A3(new_n636_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(G36gat), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n655_), .A2(KEYINPUT107), .A3(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(KEYINPUT107), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(KEYINPUT107), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n655_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n657_), .A2(new_n660_), .ZN(G1329gat));
  INV_X1    g460(.A(G43gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n642_), .B2(new_n276_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n635_), .A2(G43gat), .A3(new_n277_), .A4(new_n636_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g467(.A(G50gat), .B1(new_n646_), .B2(new_n619_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n619_), .A2(G50gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n637_), .B2(new_n670_), .ZN(G1331gat));
  INV_X1    g470(.A(G57gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n593_), .A2(new_n630_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n673_), .A2(KEYINPUT109), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n445_), .A2(new_n552_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(KEYINPUT109), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n677_), .B2(new_n440_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT110), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n538_), .A2(new_n586_), .A3(new_n630_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n680_), .A2(new_n672_), .A3(new_n440_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1332gat));
  OAI21_X1  g481(.A(G64gat), .B1(new_n680_), .B2(new_n442_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT48), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n442_), .A2(G64gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n677_), .B2(new_n685_), .ZN(G1333gat));
  OAI21_X1  g485(.A(G71gat), .B1(new_n680_), .B2(new_n276_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT49), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n276_), .A2(G71gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n677_), .B2(new_n689_), .ZN(G1334gat));
  OAI21_X1  g489(.A(G78gat), .B1(new_n680_), .B2(new_n388_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT50), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n388_), .A2(G78gat), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT111), .Z(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n677_), .B2(new_n694_), .ZN(G1335gat));
  INV_X1    g494(.A(KEYINPUT113), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n626_), .A2(KEYINPUT112), .A3(new_n628_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n582_), .A2(new_n552_), .A3(new_n631_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT112), .B1(new_n626_), .B2(new_n628_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n629_), .A2(new_n702_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n703_), .A2(KEYINPUT113), .A3(new_n698_), .A4(new_n697_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n701_), .A2(new_n411_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G85gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n640_), .A2(new_n582_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n675_), .A2(new_n707_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n440_), .A2(G85gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n708_), .B2(new_n709_), .ZN(G1336gat));
  NAND4_X1  g509(.A1(new_n701_), .A2(new_n704_), .A3(G92gat), .A4(new_n653_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n448_), .B1(new_n708_), .B2(new_n442_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT114), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1337gat));
  NAND3_X1  g513(.A1(new_n701_), .A2(new_n277_), .A3(new_n704_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G99gat), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n675_), .A2(new_n459_), .A3(new_n277_), .A4(new_n707_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT115), .Z(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT116), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n716_), .B(new_n718_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1338gat));
  AND2_X1   g524(.A1(new_n698_), .A2(new_n619_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n460_), .B1(new_n629_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n675_), .A2(new_n460_), .A3(new_n619_), .A4(new_n707_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g531(.A1(new_n552_), .A2(new_n572_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT118), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n563_), .B2(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n553_), .A2(KEYINPUT68), .A3(new_n554_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n564_), .A2(KEYINPUT12), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n481_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n740_), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(new_n557_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n739_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n554_), .B1(new_n743_), .B2(new_n553_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n558_), .B1(new_n562_), .B2(new_n561_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n557_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n735_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n744_), .B1(new_n747_), .B2(KEYINPUT117), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n563_), .A2(new_n749_), .A3(new_n735_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n742_), .A2(new_n748_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n570_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n753_), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n570_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n753_), .B1(new_n752_), .B2(new_n755_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n733_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n544_), .A2(new_n545_), .A3(new_n541_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n551_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n548_), .A2(new_n551_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n578_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n760_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n504_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT57), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n763_), .A2(new_n572_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n570_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n570_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(KEYINPUT58), .B(new_n768_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n592_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n764_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n563_), .A2(new_n749_), .A3(new_n735_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n749_), .B1(new_n563_), .B2(new_n735_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n744_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n571_), .B1(new_n779_), .B2(new_n742_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT120), .B1(new_n780_), .B2(new_n754_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n757_), .A3(new_n756_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n776_), .B1(new_n782_), .B2(new_n733_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n766_), .A2(KEYINPUT57), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n775_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n537_), .B1(new_n767_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n593_), .A2(new_n586_), .A3(new_n582_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT54), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n442_), .A2(new_n277_), .A3(new_n411_), .A4(new_n388_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n789_), .A2(KEYINPUT59), .A3(new_n791_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n586_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(G113gat), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n552_), .A2(new_n797_), .ZN(new_n798_));
  OAI22_X1  g597(.A1(new_n796_), .A2(new_n797_), .B1(new_n792_), .B2(new_n798_), .ZN(G1340gat));
  AOI21_X1  g598(.A(new_n582_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n800_));
  INV_X1    g599(.A(G120gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n582_), .B2(KEYINPUT60), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(KEYINPUT60), .B2(new_n801_), .ZN(new_n803_));
  OAI22_X1  g602(.A1(new_n800_), .A2(new_n801_), .B1(new_n792_), .B2(new_n803_), .ZN(G1341gat));
  AOI21_X1  g603(.A(new_n537_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n805_));
  INV_X1    g604(.A(G127gat), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n631_), .A2(new_n806_), .ZN(new_n807_));
  OAI22_X1  g606(.A1(new_n805_), .A2(new_n806_), .B1(new_n792_), .B2(new_n807_), .ZN(G1342gat));
  NAND2_X1  g607(.A1(new_n794_), .A2(new_n795_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n592_), .A2(G134gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT121), .ZN(new_n811_));
  INV_X1    g610(.A(G134gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n789_), .A2(new_n504_), .A3(new_n791_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n809_), .A2(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(G1343gat));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n787_), .B(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n783_), .B2(new_n504_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n504_), .A2(new_n817_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n765_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n820_), .A3(new_n775_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n816_), .B1(new_n821_), .B2(new_n537_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n277_), .A2(new_n388_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n653_), .A2(new_n440_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n356_), .A3(new_n552_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G141gat), .B1(new_n827_), .B2(new_n586_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1344gat));
  NAND3_X1  g630(.A1(new_n828_), .A2(new_n357_), .A3(new_n630_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G148gat), .B1(new_n827_), .B2(new_n582_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1345gat));
  XNOR2_X1  g633(.A(KEYINPUT61), .B(G155gat), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n828_), .A2(new_n631_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n827_), .B2(new_n537_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(G1346gat));
  NAND2_X1  g638(.A1(new_n592_), .A2(G162gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT122), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n825_), .A2(new_n504_), .A3(new_n826_), .ZN(new_n842_));
  INV_X1    g641(.A(G162gat), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n828_), .A2(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(G1347gat));
  XNOR2_X1  g643(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n276_), .A2(new_n619_), .A3(new_n411_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n653_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n552_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n845_), .B1(new_n850_), .B2(new_n236_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n845_), .ZN(new_n852_));
  OAI211_X1 g651(.A(G169gat), .B(new_n852_), .C1(new_n822_), .C2(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n211_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT124), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n851_), .A2(new_n853_), .A3(new_n857_), .A4(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1348gat));
  NAND2_X1  g658(.A1(new_n789_), .A2(new_n848_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n212_), .A2(KEYINPUT125), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n860_), .A2(new_n582_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n860_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n630_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT125), .B(G176gat), .Z(new_n865_));
  AOI21_X1  g664(.A(new_n862_), .B1(new_n864_), .B2(new_n865_), .ZN(G1349gat));
  AOI21_X1  g665(.A(G183gat), .B1(new_n863_), .B2(new_n631_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n860_), .A2(new_n228_), .A3(new_n537_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1350gat));
  AOI21_X1  g668(.A(new_n860_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n504_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n871_));
  OAI22_X1  g670(.A1(new_n870_), .A2(new_n220_), .B1(new_n860_), .B2(new_n871_), .ZN(G1351gat));
  NOR2_X1   g671(.A1(new_n442_), .A2(new_n411_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI211_X1 g673(.A(new_n824_), .B(new_n874_), .C1(new_n786_), .C2(new_n788_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n552_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g676(.A1(new_n789_), .A2(new_n823_), .A3(new_n873_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n878_), .A2(new_n582_), .A3(new_n284_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G204gat), .B1(new_n875_), .B2(new_n630_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1353gat));
  AOI211_X1 g680(.A(KEYINPUT63), .B(G211gat), .C1(new_n875_), .C2(new_n631_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT63), .B(G211gat), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n878_), .A2(new_n537_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1354gat));
  XOR2_X1   g684(.A(KEYINPUT126), .B(G218gat), .Z(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n875_), .B2(new_n504_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n592_), .A2(new_n886_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n878_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT127), .B1(new_n887_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n888_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n875_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n893_));
  NOR4_X1   g692(.A1(new_n822_), .A2(new_n766_), .A3(new_n824_), .A4(new_n874_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n892_), .B(new_n893_), .C1(new_n894_), .C2(new_n886_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n890_), .A2(new_n895_), .ZN(G1355gat));
endmodule


