//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n974_, new_n975_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n984_, new_n985_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n996_, new_n997_, new_n998_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT30), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  INV_X1    g004(.A(G15gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT25), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT77), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G183gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n210_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n209_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n222_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT77), .B(G183gat), .ZN(new_n231_));
  INV_X1    g030(.A(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n227_), .A2(new_n228_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G169gat), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n217_), .A2(new_n230_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n208_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n208_), .A2(new_n238_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT31), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT31), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n239_), .A2(new_n240_), .A3(new_n244_), .A4(new_n241_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n247_), .A2(new_n248_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n247_), .A2(new_n248_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n243_), .A2(new_n253_), .A3(new_n245_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G1gat), .B(G29gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT89), .B(KEYINPUT0), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G57gat), .B(G85gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262_));
  INV_X1    g061(.A(G141gat), .ZN(new_n263_));
  INV_X1    g062(.A(G148gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n265_), .A2(new_n268_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n263_), .A2(new_n264_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n266_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n272_), .A2(new_n279_), .A3(new_n273_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n253_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n271_), .A2(new_n274_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n249_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G225gat), .A2(G233gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT88), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT87), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(new_n283_), .B2(KEYINPUT4), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n283_), .A2(new_n285_), .A3(KEYINPUT4), .ZN(new_n291_));
  INV_X1    g090(.A(new_n287_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n282_), .A2(new_n253_), .A3(KEYINPUT87), .A4(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .A4(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n288_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT88), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n261_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n284_), .A2(new_n249_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT87), .B1(new_n300_), .B2(new_n293_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n294_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(KEYINPUT88), .A3(new_n292_), .A4(new_n291_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n288_), .A2(new_n295_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n260_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n284_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT79), .B(KEYINPUT28), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G22gat), .B(G50gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n309_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G78gat), .B(G106gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT21), .ZN(new_n316_));
  INV_X1    g115(.A(G197gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT80), .ZN(new_n318_));
  INV_X1    g117(.A(G204gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(KEYINPUT80), .A2(G204gat), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n317_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G197gat), .A2(G204gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n316_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G218gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G211gat), .ZN(new_n326_));
  INV_X1    g125(.A(G211gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G218gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n320_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n316_), .B1(G197gat), .B2(G204gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n320_), .A2(new_n321_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n323_), .B1(new_n333_), .B2(G197gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n316_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n324_), .A2(new_n332_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n308_), .B1(new_n275_), .B2(new_n281_), .ZN(new_n337_));
  OAI211_X1 g136(.A(G228gat), .B(G233gat), .C1(new_n336_), .C2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n324_), .A2(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n335_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n282_), .A2(KEYINPUT29), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G228gat), .A2(G233gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n315_), .B1(new_n338_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n313_), .B1(new_n345_), .B2(KEYINPUT81), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n338_), .A2(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n314_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n338_), .A2(new_n344_), .A3(new_n315_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n348_), .A2(KEYINPUT81), .A3(new_n349_), .A4(new_n313_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n211_), .A2(new_n232_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n227_), .A2(new_n228_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT83), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n227_), .A2(new_n354_), .A3(KEYINPUT83), .A4(new_n228_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n237_), .A3(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT25), .B(G183gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n209_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n221_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n361_), .A2(new_n234_), .A3(new_n362_), .A4(new_n224_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n341_), .A2(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n212_), .A2(new_n214_), .A3(new_n232_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n227_), .A2(new_n228_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n237_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n230_), .A2(new_n217_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n336_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n370_), .A3(KEYINPUT20), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT20), .B(new_n374_), .C1(new_n238_), .C2(new_n336_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n339_), .A2(new_n359_), .A3(new_n340_), .A4(new_n363_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT84), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  INV_X1    g180(.A(new_n209_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n213_), .A2(G183gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n211_), .A2(KEYINPUT77), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT25), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n216_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n382_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n234_), .A2(new_n362_), .A3(new_n224_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n368_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n381_), .B1(new_n341_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n378_), .A4(new_n374_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n376_), .A2(new_n380_), .A3(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n394_), .A2(KEYINPUT86), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(KEYINPUT86), .ZN(new_n396_));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397_));
  OR3_X1    g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n394_), .B(KEYINPUT86), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n397_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n399_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n393_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n376_), .A2(new_n380_), .A3(new_n392_), .A4(new_n404_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n407_), .A2(KEYINPUT27), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n365_), .A2(new_n370_), .A3(KEYINPUT20), .A4(new_n374_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT92), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n381_), .B1(new_n238_), .B2(new_n336_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n374_), .A4(new_n365_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT20), .B1(new_n238_), .B2(new_n336_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n341_), .B1(KEYINPUT91), .B2(new_n364_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n364_), .A2(KEYINPUT91), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n413_), .B(new_n416_), .C1(new_n420_), .C2(new_n374_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n405_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n411_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n410_), .A2(new_n423_), .ZN(new_n424_));
  NOR4_X1   g223(.A1(new_n255_), .A2(new_n307_), .A3(new_n353_), .A4(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT94), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT93), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n421_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n427_), .B1(new_n421_), .B2(new_n428_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n393_), .A2(new_n428_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n299_), .B2(new_n306_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n299_), .A2(KEYINPUT33), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n304_), .A2(new_n305_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n261_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n287_), .B1(new_n286_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n440_), .B2(new_n286_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n303_), .A2(new_n287_), .A3(new_n291_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n260_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n406_), .A2(new_n444_), .A3(new_n407_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n432_), .A2(new_n434_), .B1(new_n439_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n426_), .B1(new_n446_), .B2(new_n353_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT96), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n353_), .A2(new_n299_), .A3(new_n306_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n424_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n449_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n408_), .A2(new_n409_), .B1(new_n411_), .B2(new_n422_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT96), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n341_), .A2(new_n389_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n455_), .A2(KEYINPUT20), .A3(new_n378_), .A4(new_n374_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n456_), .A2(KEYINPUT84), .B1(new_n371_), .B2(new_n375_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n404_), .B1(new_n457_), .B2(new_n392_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n407_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n437_), .B1(new_n436_), .B2(new_n261_), .ZN(new_n461_));
  AOI211_X1 g260(.A(KEYINPUT33), .B(new_n260_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n460_), .B(new_n444_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n421_), .A2(new_n428_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT93), .ZN(new_n465_));
  INV_X1    g264(.A(new_n433_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n307_), .A3(new_n466_), .A4(new_n429_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n353_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT94), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n447_), .A2(new_n454_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n425_), .B1(new_n470_), .B2(new_n255_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n474_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT75), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G1gat), .B(G8gat), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n476_), .A2(new_n477_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n479_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n480_), .A2(new_n481_), .A3(new_n490_), .A4(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n490_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n491_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n480_), .A2(new_n493_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT75), .B1(new_n499_), .B2(new_n495_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n490_), .A2(new_n478_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n498_), .B1(new_n496_), .B2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n503_), .A2(KEYINPUT74), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(KEYINPUT74), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT76), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G169gat), .B(G197gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n501_), .A2(new_n504_), .A3(new_n505_), .A4(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(G230gat), .A2(G233gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT6), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(G99gat), .A3(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(G85gat), .A3(G92gat), .ZN(new_n523_));
  INV_X1    g322(.A(G85gat), .ZN(new_n524_));
  INV_X1    g323(.A(G92gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n521_), .B(new_n523_), .C1(new_n528_), .C2(new_n522_), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT10), .B(G99gat), .Z(new_n530_));
  INV_X1    g329(.A(G106gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(KEYINPUT64), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT64), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT10), .B(G99gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n533_), .B1(new_n534_), .B2(G106gat), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n529_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(G99gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(new_n531_), .A3(KEYINPUT65), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT7), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT7), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n540_), .A2(new_n537_), .A3(new_n531_), .A4(KEYINPUT65), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n521_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n528_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT8), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT8), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n546_), .A3(new_n543_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n536_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G57gat), .B(G64gat), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n549_), .A2(KEYINPUT11), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(KEYINPUT11), .ZN(new_n551_));
  XOR2_X1   g350(.A(G71gat), .B(G78gat), .Z(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n551_), .A2(new_n552_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n532_), .A2(new_n535_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n543_), .A2(KEYINPUT9), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n521_), .A2(new_n523_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n546_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n542_), .A2(new_n546_), .A3(new_n543_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n560_), .B(new_n555_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n516_), .B1(new_n556_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT66), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n562_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT66), .B1(new_n545_), .B2(new_n547_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n560_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n555_), .A2(KEYINPUT67), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT67), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n553_), .A2(new_n571_), .A3(new_n554_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n570_), .A2(KEYINPUT12), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT68), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n569_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n566_), .B1(new_n562_), .B2(new_n561_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n545_), .A2(KEYINPUT66), .A3(new_n547_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n536_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n570_), .A2(KEYINPUT12), .A3(new_n572_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT68), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n560_), .B1(new_n562_), .B2(new_n561_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n555_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT12), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n564_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n575_), .A2(new_n580_), .A3(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n565_), .B1(new_n585_), .B2(new_n516_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G120gat), .B(G148gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(KEYINPUT13), .A3(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n471_), .A2(new_n515_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT34), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT35), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n576_), .A2(new_n577_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n499_), .B1(new_n604_), .B2(new_n560_), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n581_), .A2(new_n478_), .B1(KEYINPUT35), .B2(new_n601_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n601_), .A2(KEYINPUT35), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n548_), .B2(new_n491_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n609_), .B(new_n602_), .C1(new_n499_), .C2(new_n578_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G134gat), .B(G162gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT70), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n607_), .A2(new_n610_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n607_), .A2(new_n610_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n613_), .B(KEYINPUT36), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n617_), .A2(KEYINPUT71), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT71), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n607_), .A2(new_n621_), .A3(new_n610_), .A4(new_n616_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n599_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n619_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n617_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n623_), .A2(KEYINPUT73), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT73), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n617_), .A2(KEYINPUT71), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n624_), .A3(new_n622_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT37), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n629_), .B1(new_n632_), .B2(new_n626_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n628_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n582_), .A2(new_n490_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n495_), .A2(new_n555_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(G231gat), .ZN(new_n638_));
  INV_X1    g437(.A(G233gat), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n635_), .A2(new_n636_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(G127gat), .B(G155gat), .Z(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT16), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G183gat), .B(G211gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT17), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n647_), .A2(new_n571_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n643_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n648_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n634_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n598_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n483_), .A3(new_n307_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT38), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n624_), .A2(new_n617_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(KEYINPUT97), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(KEYINPUT97), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n655_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n598_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n307_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G1gat), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n659_), .A2(new_n668_), .ZN(G1324gat));
  NAND3_X1  g468(.A1(new_n657_), .A2(new_n484_), .A3(new_n424_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n598_), .A2(new_n424_), .A3(new_n664_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G8gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT98), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n675_), .A3(G8gat), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n673_), .A2(new_n674_), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n674_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n670_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT40), .B(new_n670_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1325gat));
  INV_X1    g482(.A(new_n255_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n657_), .A2(new_n206_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n665_), .A2(new_n684_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n686_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT41), .B1(new_n686_), .B2(G15gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1326gat));
  INV_X1    g490(.A(G22gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n665_), .B2(new_n353_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT42), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n657_), .A2(new_n692_), .A3(new_n353_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1327gat));
  INV_X1    g495(.A(new_n663_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n654_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n598_), .A2(new_n698_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n699_), .A2(G29gat), .A3(new_n667_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n451_), .A2(new_n452_), .A3(KEYINPUT96), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n448_), .B1(new_n424_), .B2(new_n449_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n703_), .B(new_n704_), .C1(new_n468_), .C2(KEYINPUT94), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n446_), .A2(new_n426_), .A3(new_n353_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n255_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n425_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n702_), .B1(new_n709_), .B2(new_n634_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT73), .B1(new_n623_), .B2(new_n627_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n632_), .A2(new_n629_), .A3(new_n626_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AOI211_X1 g512(.A(KEYINPUT43), .B(new_n713_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n710_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n597_), .A2(new_n515_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n655_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n701_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n471_), .B2(new_n713_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n463_), .A2(new_n467_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n353_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT94), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n704_), .A2(new_n703_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n684_), .B1(new_n724_), .B2(new_n469_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n702_), .B(new_n634_), .C1(new_n725_), .C2(new_n425_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n719_), .A2(new_n726_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n727_), .A2(KEYINPUT44), .A3(new_n716_), .A4(new_n655_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n718_), .A2(new_n307_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n700_), .B1(new_n729_), .B2(G29gat), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT100), .ZN(G1328gat));
  XNOR2_X1  g530(.A(new_n424_), .B(KEYINPUT101), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(G36gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n598_), .A2(new_n698_), .A3(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT45), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n718_), .A2(new_n424_), .A3(new_n728_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(G36gat), .B2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n737_), .B(new_n739_), .ZN(G1329gat));
  AND4_X1   g539(.A1(G43gat), .A2(new_n718_), .A3(new_n684_), .A4(new_n728_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n699_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G43gat), .B1(new_n742_), .B2(new_n684_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(G1330gat));
  NOR3_X1   g545(.A1(new_n699_), .A2(G50gat), .A3(new_n721_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n718_), .A2(new_n353_), .A3(new_n728_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G50gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT104), .ZN(G1331gat));
  INV_X1    g549(.A(new_n597_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n471_), .A2(new_n514_), .A3(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(new_n664_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G57gat), .B1(new_n754_), .B2(new_n667_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n752_), .A2(new_n656_), .ZN(new_n756_));
  INV_X1    g555(.A(G57gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n307_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1332gat));
  INV_X1    g558(.A(G64gat), .ZN(new_n760_));
  INV_X1    g559(.A(new_n732_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n753_), .A2(new_n761_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G64gat), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(KEYINPUT48), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(KEYINPUT48), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT105), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(new_n762_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n753_), .B2(new_n684_), .ZN(new_n773_));
  XOR2_X1   g572(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n756_), .A2(new_n772_), .A3(new_n684_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1334gat));
  INV_X1    g576(.A(G78gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n753_), .B2(new_n353_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT50), .Z(new_n780_));
  NAND2_X1  g579(.A1(new_n353_), .A2(new_n778_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT107), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n756_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(G1335gat));
  NOR3_X1   g583(.A1(new_n751_), .A2(new_n514_), .A3(new_n654_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n727_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n667_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n752_), .A2(new_n698_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n307_), .A2(new_n524_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT108), .ZN(G1336gat));
  OAI21_X1  g590(.A(G92gat), .B1(new_n786_), .B2(new_n732_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n788_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n525_), .A3(new_n424_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1337gat));
  OAI21_X1  g594(.A(G99gat), .B1(new_n786_), .B2(new_n255_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n752_), .A2(new_n530_), .A3(new_n684_), .A4(new_n698_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT109), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT111), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(KEYINPUT110), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n798_), .B(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n796_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n800_), .A2(new_n802_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n802_), .B1(new_n800_), .B2(new_n806_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n793_), .A2(new_n531_), .A3(new_n353_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n353_), .B(new_n785_), .C1(new_n710_), .C2(new_n714_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(G106gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(G106gat), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n813_), .A2(new_n814_), .A3(KEYINPUT52), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  INV_X1    g615(.A(new_n785_), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n721_), .B(new_n817_), .C1(new_n719_), .C2(new_n726_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT112), .B1(new_n818_), .B2(new_n531_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n811_), .A2(new_n812_), .A3(G106gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n810_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT53), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n810_), .C1(new_n815_), .C2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1339gat));
  NAND2_X1  g625(.A1(new_n591_), .A2(new_n514_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n516_), .A2(KEYINPUT114), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n575_), .A2(new_n580_), .A3(new_n584_), .A4(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n585_), .B2(new_n828_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n585_), .A2(new_n516_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n590_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n590_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n827_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n496_), .A2(new_n502_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n510_), .B1(new_n840_), .B2(new_n498_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n497_), .A2(new_n500_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n498_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n513_), .A2(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n593_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n697_), .B1(new_n839_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n591_), .A2(new_n844_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n590_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT56), .B1(new_n834_), .B2(new_n590_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT58), .B(new_n849_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(KEYINPUT115), .A3(new_n634_), .A4(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n697_), .B(KEYINPUT57), .C1(new_n839_), .C2(new_n845_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n848_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n713_), .B1(new_n853_), .B2(new_n852_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT115), .B1(new_n859_), .B2(new_n855_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n655_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n654_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n864_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n713_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n865_), .B2(new_n713_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n861_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n861_), .A2(KEYINPUT116), .A3(new_n870_), .ZN(new_n874_));
  NOR4_X1   g673(.A1(new_n255_), .A2(new_n667_), .A3(new_n353_), .A4(new_n424_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n514_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n854_), .A2(new_n634_), .A3(new_n855_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n848_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n848_), .A2(KEYINPUT117), .A3(new_n879_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(new_n857_), .A3(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n869_), .B1(new_n884_), .B2(new_n655_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n875_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n879_), .A2(new_n889_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n890_), .A2(new_n856_), .A3(new_n848_), .A4(new_n857_), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n872_), .B(new_n869_), .C1(new_n891_), .C2(new_n655_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT116), .B1(new_n861_), .B2(new_n870_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n875_), .ZN(new_n895_));
  AOI211_X1 g694(.A(new_n515_), .B(new_n888_), .C1(new_n895_), .C2(KEYINPUT59), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n878_), .B1(new_n896_), .B2(new_n877_), .ZN(G1340gat));
  AOI211_X1 g696(.A(new_n751_), .B(new_n888_), .C1(new_n895_), .C2(KEYINPUT59), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT118), .B(G120gat), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(KEYINPUT60), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n751_), .A2(KEYINPUT60), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n899_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n876_), .B2(new_n903_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n876_), .A2(new_n900_), .A3(new_n903_), .ZN(new_n905_));
  OAI22_X1  g704(.A1(new_n898_), .A2(new_n899_), .B1(new_n904_), .B2(new_n905_), .ZN(G1341gat));
  INV_X1    g705(.A(new_n888_), .ZN(new_n907_));
  INV_X1    g706(.A(G127gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n655_), .A2(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n907_), .B(new_n909_), .C1(new_n876_), .C2(new_n886_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n873_), .A2(new_n654_), .A3(new_n874_), .A4(new_n875_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n908_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT120), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n912_), .A2(KEYINPUT120), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1342gat));
  AOI21_X1  g715(.A(G134gat), .B1(new_n876_), .B2(new_n663_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n888_), .B1(new_n895_), .B2(KEYINPUT59), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n634_), .A2(G134gat), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT121), .Z(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n918_), .B2(new_n920_), .ZN(G1343gat));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n684_), .A2(new_n721_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n924_), .A2(new_n667_), .A3(new_n761_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n922_), .B1(new_n894_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n892_), .A2(new_n893_), .A3(KEYINPUT122), .A4(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n514_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT123), .B(G141gat), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n514_), .B(new_n930_), .C1(new_n926_), .C2(new_n928_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1344gat));
  OAI21_X1  g733(.A(new_n597_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(G148gat), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n264_), .B(new_n597_), .C1(new_n926_), .C2(new_n928_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1345gat));
  OAI21_X1  g737(.A(new_n654_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n940_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n654_), .B(new_n942_), .C1(new_n926_), .C2(new_n928_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1346gat));
  INV_X1    g743(.A(G162gat), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n945_), .B(new_n663_), .C1(new_n926_), .C2(new_n928_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n873_), .A2(new_n874_), .ZN(new_n947_));
  OAI21_X1  g746(.A(KEYINPUT122), .B1(new_n947_), .B2(new_n927_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n894_), .A2(new_n922_), .A3(new_n925_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n713_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n946_), .B1(new_n950_), .B2(new_n945_), .ZN(G1347gat));
  NAND2_X1  g750(.A1(new_n884_), .A2(new_n655_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n870_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n732_), .A2(new_n307_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n684_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n955_), .A2(new_n353_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n953_), .A2(new_n514_), .A3(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT62), .B1(new_n957_), .B2(KEYINPUT22), .ZN(new_n958_));
  OAI21_X1  g757(.A(G169gat), .B1(new_n957_), .B2(KEYINPUT62), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n960_), .B1(new_n218_), .B2(new_n958_), .ZN(G1348gat));
  NOR3_X1   g760(.A1(new_n885_), .A2(new_n353_), .A3(new_n955_), .ZN(new_n962_));
  AOI21_X1  g761(.A(G176gat), .B1(new_n962_), .B2(new_n597_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n947_), .A2(new_n353_), .ZN(new_n964_));
  NOR3_X1   g763(.A1(new_n955_), .A2(new_n219_), .A3(new_n751_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n964_), .B2(new_n965_), .ZN(G1349gat));
  NOR2_X1   g765(.A1(new_n655_), .A2(new_n360_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n953_), .A2(new_n956_), .A3(new_n967_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(KEYINPUT124), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n955_), .A2(new_n655_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n964_), .A2(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n971_), .A2(new_n231_), .ZN(new_n972_));
  AND2_X1   g771(.A1(new_n969_), .A2(new_n972_), .ZN(G1350gat));
  NAND3_X1  g772(.A1(new_n962_), .A2(new_n209_), .A3(new_n663_), .ZN(new_n974_));
  AND2_X1   g773(.A1(new_n962_), .A2(new_n634_), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n974_), .B1(new_n975_), .B2(new_n232_), .ZN(G1351gat));
  INV_X1    g775(.A(new_n954_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n924_), .A2(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(new_n978_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n947_), .A2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n980_), .A2(new_n514_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(KEYINPUT125), .B(G197gat), .ZN(new_n982_));
  XNOR2_X1  g781(.A(new_n981_), .B(new_n982_), .ZN(G1352gat));
  NOR3_X1   g782(.A1(new_n947_), .A2(new_n751_), .A3(new_n979_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n984_), .A2(G204gat), .ZN(new_n985_));
  AOI21_X1  g784(.A(new_n985_), .B1(new_n333_), .B2(new_n984_), .ZN(G1353gat));
  NAND3_X1  g785(.A1(new_n894_), .A2(new_n654_), .A3(new_n978_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n988_));
  AND2_X1   g787(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n989_));
  NOR3_X1   g788(.A1(new_n987_), .A2(new_n988_), .A3(new_n989_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n987_), .A2(new_n988_), .ZN(new_n991_));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n991_), .A2(new_n992_), .ZN(new_n993_));
  NAND3_X1  g792(.A1(new_n987_), .A2(KEYINPUT126), .A3(new_n988_), .ZN(new_n994_));
  AOI21_X1  g793(.A(new_n990_), .B1(new_n993_), .B2(new_n994_), .ZN(G1354gat));
  AOI21_X1  g794(.A(G218gat), .B1(new_n980_), .B2(new_n663_), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n634_), .A2(G218gat), .ZN(new_n997_));
  XNOR2_X1  g796(.A(new_n997_), .B(KEYINPUT127), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n996_), .B1(new_n980_), .B2(new_n998_), .ZN(G1355gat));
endmodule


