//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n206_), .B(KEYINPUT71), .ZN(new_n211_));
  INV_X1    g010(.A(new_n209_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G29gat), .B(G36gat), .Z(new_n215_));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT15), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n220_), .B(new_n221_), .C1(new_n214_), .C2(new_n217_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n214_), .B(new_n217_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT72), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n222_), .B1(new_n225_), .B2(new_n221_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G141gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G197gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n227_), .B(new_n228_), .Z(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n226_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n222_), .B(new_n229_), .C1(new_n225_), .C2(new_n221_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G230gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  AND3_X1   g036(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G99gat), .ZN(new_n241_));
  INV_X1    g040(.A(G106gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT66), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT7), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT7), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n245_), .A2(new_n241_), .A3(new_n242_), .A4(KEYINPUT66), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n240_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G85gat), .B(G92gat), .Z(new_n248_));
  AOI21_X1  g047(.A(new_n237_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n237_), .A3(new_n248_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n240_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT65), .B(G85gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G92gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT64), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n263_), .A3(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n242_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n250_), .A2(new_n251_), .B1(new_n258_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G57gat), .B(G64gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT11), .ZN(new_n269_));
  XOR2_X1   g068(.A(G71gat), .B(G78gat), .Z(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n268_), .A2(KEYINPUT11), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n269_), .A2(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n267_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n267_), .A2(new_n275_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n236_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT12), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n267_), .B2(new_n275_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n251_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT67), .B1(new_n282_), .B2(new_n249_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n250_), .A2(new_n284_), .A3(new_n251_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n283_), .A2(new_n285_), .B1(new_n266_), .B2(new_n258_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n273_), .A2(KEYINPUT12), .A3(new_n274_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n281_), .B(new_n276_), .C1(new_n286_), .C2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n279_), .B1(new_n288_), .B2(new_n236_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G120gat), .B(G148gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G176gat), .B(G204gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n289_), .B(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n295_), .A2(KEYINPUT13), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(KEYINPUT13), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n234_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  INV_X1    g105(.A(G155gat), .ZN(new_n307_));
  INV_X1    g106(.A(G162gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n306_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT1), .B1(new_n307_), .B2(new_n308_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n305_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n302_), .A2(new_n317_), .B1(new_n304_), .B2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n316_), .B(new_n319_), .C1(new_n318_), .C2(new_n304_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n309_), .A2(new_n306_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n313_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT28), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G22gat), .B(G50gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n325_), .B(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT80), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n325_), .B(new_n326_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G211gat), .B(G218gat), .ZN(new_n333_));
  INV_X1    g132(.A(G197gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G204gat), .ZN(new_n335_));
  INV_X1    g134(.A(G204gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G197gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(KEYINPUT81), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT81), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT21), .B1(new_n335_), .B2(new_n340_), .ZN(new_n341_));
  OAI221_X1 g140(.A(new_n333_), .B1(KEYINPUT21), .B2(new_n338_), .C1(new_n339_), .C2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n333_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(KEYINPUT21), .A3(new_n338_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n346_));
  AND2_X1   g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n346_), .A2(new_n347_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G78gat), .B(G106gat), .Z(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT82), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OR3_X1    g151(.A1(new_n348_), .A2(new_n349_), .A3(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n352_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n329_), .A2(new_n332_), .A3(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n354_), .A2(KEYINPUT83), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(KEYINPUT83), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n357_), .A2(new_n330_), .A3(new_n353_), .A4(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT20), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366_));
  INV_X1    g165(.A(G169gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT22), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT22), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G169gat), .ZN(new_n370_));
  INV_X1    g169(.A(G176gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G183gat), .ZN(new_n373_));
  INV_X1    g172(.A(G190gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT23), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT74), .B(KEYINPUT23), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n376_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n366_), .B(new_n372_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n366_), .ZN(new_n385_));
  MUX2_X1   g184(.A(new_n384_), .B(new_n385_), .S(KEYINPUT24), .Z(new_n386_));
  NAND2_X1  g185(.A1(new_n375_), .A2(new_n377_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n379_), .B2(new_n375_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT73), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT26), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(G190gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT26), .B(G190gat), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n389_), .B(new_n392_), .C1(new_n393_), .C2(new_n390_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n386_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n382_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n365_), .B1(new_n396_), .B2(new_n345_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n383_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n385_), .B2(new_n398_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n380_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n389_), .B(KEYINPUT86), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n402_), .A2(new_n393_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT89), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n369_), .A2(G169gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n367_), .A2(KEYINPUT22), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n368_), .A2(new_n370_), .A3(KEYINPUT89), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n371_), .A3(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n366_), .B(KEYINPUT88), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT90), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT90), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n381_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n388_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n406_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n412_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n416_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n406_), .B(new_n420_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n405_), .B1(new_n421_), .B2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n364_), .B(new_n397_), .C1(new_n426_), .C2(new_n345_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n345_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n395_), .A3(new_n382_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT20), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(KEYINPUT92), .A3(new_n345_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT92), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT91), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n404_), .B1(new_n434_), .B2(new_n424_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n432_), .B1(new_n435_), .B2(new_n428_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n430_), .B1(new_n431_), .B2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n363_), .B(KEYINPUT85), .Z(new_n438_));
  OAI21_X1  g237(.A(new_n427_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G8gat), .B(G36gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(G64gat), .B(G92gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n439_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n444_), .B(new_n427_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT27), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n430_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT92), .B1(new_n426_), .B2(new_n345_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n435_), .A2(new_n432_), .A3(new_n428_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n451_), .B(new_n438_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT96), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT96), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n437_), .A2(new_n456_), .A3(new_n438_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n405_), .A2(new_n428_), .A3(new_n433_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n364_), .B1(new_n458_), .B2(new_n397_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n455_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT97), .A3(new_n445_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n447_), .A2(KEYINPUT27), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n459_), .B1(new_n454_), .B2(KEYINPUT96), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n444_), .B1(new_n466_), .B2(new_n457_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(KEYINPUT97), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n360_), .B(new_n450_), .C1(new_n465_), .C2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT98), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT4), .ZN(new_n473_));
  XOR2_X1   g272(.A(G127gat), .B(G134gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(G113gat), .B(G120gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n322_), .A2(KEYINPUT94), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n476_), .B(new_n477_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(KEYINPUT94), .A3(new_n322_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n473_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n478_), .A2(new_n322_), .A3(KEYINPUT4), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n472_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n480_), .A2(new_n482_), .A3(new_n471_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G1gat), .B(G29gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(G85gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT0), .B(G57gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n487_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n463_), .B1(new_n467_), .B2(KEYINPUT97), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n461_), .A2(new_n445_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT98), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n360_), .A4(new_n450_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G15gat), .B(G43gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT75), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT30), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(new_n396_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(new_n478_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G227gat), .A2(G233gat), .ZN(new_n506_));
  INV_X1    g305(.A(G71gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(new_n241_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT31), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n505_), .B(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n470_), .A2(new_n493_), .A3(new_n500_), .A4(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n360_), .A2(new_n492_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n513_), .B(new_n450_), .C1(new_n465_), .C2(new_n468_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n491_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n516_), .A2(KEYINPUT33), .ZN(new_n517_));
  OR3_X1    g316(.A1(new_n483_), .A2(new_n472_), .A3(new_n484_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n480_), .A2(new_n482_), .A3(KEYINPUT95), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT95), .B1(new_n480_), .B2(new_n482_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n472_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n515_), .A3(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n516_), .B2(KEYINPUT33), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n448_), .A2(new_n517_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n444_), .A2(KEYINPUT32), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n487_), .A2(new_n491_), .ZN(new_n527_));
  OAI22_X1  g326(.A1(new_n439_), .A2(new_n526_), .B1(new_n527_), .B2(new_n516_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n526_), .B2(new_n461_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n360_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n514_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n511_), .B(KEYINPUT78), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n301_), .B1(new_n512_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n267_), .ZN(new_n535_));
  OAI22_X1  g334(.A1(new_n286_), .A2(new_n218_), .B1(new_n217_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n542_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G134gat), .B(G162gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n536_), .A2(new_n545_), .B1(KEYINPUT36), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n548_), .A2(KEYINPUT36), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n275_), .B(new_n557_), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(new_n214_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561_));
  XOR2_X1   g360(.A(G127gat), .B(G155gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT16), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n560_), .A2(new_n561_), .A3(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(KEYINPUT17), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n560_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n556_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n534_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(new_n202_), .A3(new_n492_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT38), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n554_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n512_), .B2(new_n533_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n301_), .A2(new_n569_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G1gat), .B1(new_n579_), .B2(new_n493_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n572_), .A2(new_n573_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n574_), .A2(new_n580_), .A3(new_n581_), .ZN(G1324gat));
  NAND2_X1  g381(.A1(new_n498_), .A2(new_n450_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n571_), .A2(new_n203_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n583_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G8gat), .B1(new_n579_), .B2(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n586_), .A2(KEYINPUT39), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(KEYINPUT39), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n584_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g389(.A(G15gat), .ZN(new_n591_));
  INV_X1    g390(.A(new_n532_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n578_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT99), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT41), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n571_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT100), .Z(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n597_), .A3(new_n599_), .ZN(G1326gat));
  INV_X1    g399(.A(G22gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n360_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n571_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G22gat), .B1(new_n579_), .B2(new_n360_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(KEYINPUT42), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(KEYINPUT42), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT101), .Z(G1327gat));
  INV_X1    g407(.A(new_n569_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n554_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n534_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(G29gat), .B1(new_n611_), .B2(new_n492_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n301_), .A2(new_n609_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n512_), .A2(new_n533_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n615_), .B2(new_n556_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n556_), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT43), .B(new_n617_), .C1(new_n512_), .C2(new_n533_), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT44), .B(new_n613_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n619_), .A2(G29gat), .A3(new_n492_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n613_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n612_), .B1(new_n620_), .B2(new_n623_), .ZN(G1328gat));
  INV_X1    g423(.A(G36gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n611_), .A2(new_n625_), .A3(new_n583_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT45), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n617_), .B1(new_n512_), .B2(new_n533_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(new_n614_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT44), .B1(new_n630_), .B2(new_n613_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n619_), .A2(new_n583_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n628_), .B(G36gat), .C1(new_n631_), .C2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n623_), .A2(new_n583_), .A3(new_n619_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n628_), .B1(new_n635_), .B2(G36gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n627_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI221_X1 g438(.A(new_n627_), .B1(KEYINPUT103), .B2(KEYINPUT46), .C1(new_n634_), .C2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1329gat));
  XOR2_X1   g440(.A(KEYINPUT104), .B(G43gat), .Z(new_n642_));
  INV_X1    g441(.A(new_n611_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n642_), .B1(new_n643_), .B2(new_n532_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n619_), .A2(G43gat), .A3(new_n511_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(new_n631_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(G1330gat));
  NAND2_X1  g447(.A1(new_n619_), .A2(new_n602_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G50gat), .B1(new_n631_), .B2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n360_), .A2(G50gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT106), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n643_), .B2(new_n652_), .ZN(G1331gat));
  AOI211_X1 g452(.A(new_n233_), .B(new_n298_), .C1(new_n512_), .C2(new_n533_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n570_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT107), .Z(new_n656_));
  AOI21_X1  g455(.A(G57gat), .B1(new_n656_), .B2(new_n492_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n233_), .A2(new_n569_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n576_), .A2(new_n299_), .A3(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(G57gat), .A3(new_n492_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT108), .Z(new_n661_));
  NOR2_X1   g460(.A1(new_n657_), .A2(new_n661_), .ZN(G1332gat));
  INV_X1    g461(.A(G64gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n659_), .B2(new_n583_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT48), .Z(new_n665_));
  NAND3_X1  g464(.A1(new_n656_), .A2(new_n663_), .A3(new_n583_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1333gat));
  AOI21_X1  g466(.A(new_n507_), .B1(new_n659_), .B2(new_n592_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT49), .Z(new_n669_));
  NAND3_X1  g468(.A1(new_n656_), .A2(new_n507_), .A3(new_n592_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1334gat));
  INV_X1    g470(.A(G78gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n659_), .B2(new_n602_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT50), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n656_), .A2(new_n672_), .A3(new_n602_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1335gat));
  AND2_X1   g475(.A1(new_n654_), .A2(new_n610_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G85gat), .B1(new_n677_), .B2(new_n492_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n233_), .A2(new_n298_), .A3(new_n609_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n630_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n492_), .A2(new_n253_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1336gat));
  INV_X1    g481(.A(G92gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n677_), .A2(new_n683_), .A3(new_n583_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n680_), .A2(new_n583_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n686_), .B2(new_n683_), .ZN(G1337gat));
  AND3_X1   g486(.A1(new_n677_), .A2(new_n265_), .A3(new_n511_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n680_), .A2(new_n592_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G99gat), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g490(.A1(new_n677_), .A2(new_n242_), .A3(new_n602_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n630_), .A2(new_n602_), .A3(new_n679_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT52), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(new_n694_), .A3(G106gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n693_), .B2(G106gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT53), .ZN(G1339gat));
  OR2_X1    g497(.A1(new_n289_), .A2(new_n294_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n214_), .A2(new_n217_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n221_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n229_), .B1(new_n701_), .B2(new_n220_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n221_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n225_), .B2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n232_), .A2(new_n699_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT56), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n281_), .A2(new_n276_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n283_), .A2(new_n285_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n258_), .A2(new_n266_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n287_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n236_), .B1(new_n707_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n288_), .A2(KEYINPUT111), .A3(new_n236_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT55), .B1(new_n288_), .B2(new_n236_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n281_), .A2(new_n276_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n708_), .A2(new_n709_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n287_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT55), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n716_), .A2(new_n719_), .A3(new_n720_), .A4(new_n235_), .ZN(new_n721_));
  AOI22_X1  g520(.A1(new_n713_), .A2(new_n714_), .B1(new_n715_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n294_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n713_), .A2(new_n714_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n715_), .A2(new_n721_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n723_), .A3(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n706_), .B1(new_n724_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n726_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT112), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n722_), .A2(new_n723_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT56), .A4(new_n294_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n705_), .B1(new_n728_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n733_), .A2(new_n734_), .A3(KEYINPUT58), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT58), .B1(new_n733_), .B2(new_n734_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n556_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n724_), .B2(new_n727_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT113), .A4(new_n294_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT114), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .A4(new_n706_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n699_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n739_), .A2(new_n706_), .A3(new_n740_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n732_), .A2(KEYINPUT114), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n742_), .B(new_n744_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n232_), .A2(new_n295_), .A3(new_n704_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n575_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n737_), .B1(new_n749_), .B2(KEYINPUT57), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n751_), .B(new_n575_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n569_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n658_), .A2(KEYINPUT109), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n233_), .B2(new_n569_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(new_n298_), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT54), .B1(new_n757_), .B2(new_n556_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT110), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(KEYINPUT54), .C1(new_n757_), .C2(new_n556_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n757_), .A2(KEYINPUT54), .A3(new_n556_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n753_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n470_), .A2(new_n492_), .A3(new_n500_), .A4(new_n511_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT59), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n752_), .B1(new_n750_), .B2(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n737_), .B(KEYINPUT117), .C1(new_n749_), .C2(KEYINPUT57), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n609_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n763_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n766_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n768_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(G113gat), .B1(new_n777_), .B2(new_n234_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n234_), .A2(G113gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n767_), .B2(new_n779_), .ZN(G1340gat));
  OAI21_X1  g579(.A(G120gat), .B1(new_n777_), .B2(new_n298_), .ZN(new_n781_));
  INV_X1    g580(.A(G120gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n298_), .B2(KEYINPUT60), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(KEYINPUT60), .B2(new_n782_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n767_), .B2(new_n784_), .ZN(G1341gat));
  NAND2_X1  g584(.A1(new_n609_), .A2(G127gat), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT118), .Z(new_n787_));
  NOR2_X1   g586(.A1(new_n767_), .A2(new_n569_), .ZN(new_n788_));
  OAI22_X1  g587(.A1(new_n777_), .A2(new_n787_), .B1(G127gat), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT119), .ZN(G1342gat));
  OAI21_X1  g589(.A(G134gat), .B1(new_n777_), .B2(new_n617_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n554_), .A2(G134gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n767_), .B2(new_n792_), .ZN(G1343gat));
  AOI211_X1 g592(.A(new_n360_), .B(new_n592_), .C1(new_n753_), .C2(new_n763_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n583_), .A2(new_n493_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n234_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g597(.A1(new_n796_), .A2(new_n298_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(G148gat), .Z(G1345gat));
  XOR2_X1   g599(.A(KEYINPUT61), .B(G155gat), .Z(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n796_), .B2(new_n569_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n801_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n794_), .A2(new_n609_), .A3(new_n795_), .A4(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1346gat));
  NOR3_X1   g606(.A1(new_n796_), .A2(new_n308_), .A3(new_n617_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n308_), .B1(new_n796_), .B2(new_n554_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT122), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n810_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(G1347gat));
  NOR2_X1   g612(.A1(new_n585_), .A2(new_n492_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n592_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n602_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n233_), .B(new_n816_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n410_), .A2(new_n411_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT123), .B1(new_n817_), .B2(G169gat), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n820_), .A2(new_n821_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n817_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(G1348gat));
  AOI21_X1  g624(.A(new_n602_), .B1(new_n753_), .B2(new_n763_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n815_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n826_), .A2(G176gat), .A3(new_n299_), .A4(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n299_), .B(new_n816_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n829_), .A2(KEYINPUT124), .A3(new_n371_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT124), .B1(new_n829_), .B2(new_n371_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n828_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT125), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT125), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n828_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1349gat));
  INV_X1    g635(.A(new_n816_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n774_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n569_), .A2(new_n402_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n826_), .A2(new_n609_), .A3(new_n827_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n838_), .A2(new_n839_), .B1(new_n373_), .B2(new_n840_), .ZN(G1350gat));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n575_), .A3(new_n393_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n774_), .A2(new_n617_), .A3(new_n837_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n374_), .ZN(G1351gat));
  INV_X1    g643(.A(KEYINPUT126), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n794_), .A2(new_n814_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n233_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n848_), .B2(new_n334_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n334_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n847_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n233_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(G1352gat));
  NOR2_X1   g651(.A1(new_n846_), .A2(new_n298_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n336_), .ZN(G1353gat));
  NAND2_X1  g653(.A1(new_n847_), .A2(new_n609_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n856_));
  AND2_X1   g655(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n855_), .B2(new_n856_), .ZN(G1354gat));
  AND3_X1   g658(.A1(new_n847_), .A2(G218gat), .A3(new_n556_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT127), .B1(new_n847_), .B2(new_n575_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(G218gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n847_), .A2(KEYINPUT127), .A3(new_n575_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n862_), .B2(new_n863_), .ZN(G1355gat));
endmodule


