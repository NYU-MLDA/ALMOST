//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_;
  INV_X1    g000(.A(KEYINPUT8), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n216_));
  AND2_X1   g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n208_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n202_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n206_), .A2(new_n207_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n217_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n222_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT8), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n214_), .A2(new_n218_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(KEYINPUT9), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT64), .B(G85gat), .Z(new_n232_));
  INV_X1    g031(.A(KEYINPUT9), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(G92gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT10), .B(G99gat), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n205_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n230_), .A2(new_n231_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n223_), .A2(new_n229_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n223_), .A2(new_n229_), .A3(KEYINPUT66), .A4(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G64gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT67), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G71gat), .B(G78gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n243_), .B(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n246_), .B1(new_n250_), .B2(KEYINPUT11), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n244_), .A2(new_n245_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n248_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n252_), .A3(new_n247_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(KEYINPUT11), .A3(new_n246_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n240_), .A2(new_n259_), .A3(new_n241_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n254_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n261_), .B(new_n263_), .C1(new_n255_), .C2(new_n254_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT12), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n254_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n253_), .A2(KEYINPUT12), .A3(new_n238_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n260_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n268_), .A3(new_n262_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT5), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G176gat), .B(G204gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n264_), .A2(new_n269_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT13), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT69), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G29gat), .B(G36gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G43gat), .B(G50gat), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G15gat), .B(G22gat), .ZN(new_n287_));
  INV_X1    g086(.A(G1gat), .ZN(new_n288_));
  INV_X1    g087(.A(G8gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT14), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G1gat), .B(G8gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n286_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G229gat), .A2(G233gat), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n285_), .B(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n293_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n286_), .B(new_n293_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n295_), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n296_), .A2(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G113gat), .B(G141gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(G169gat), .B(G197gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n302_), .A2(new_n305_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n280_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT96), .B(KEYINPUT27), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G169gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(G183gat), .B2(G190gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT79), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G183gat), .A3(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n325_), .B2(new_n319_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n318_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n322_), .A2(new_n324_), .A3(KEYINPUT23), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT80), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n322_), .A2(new_n324_), .A3(KEYINPUT80), .A4(KEYINPUT23), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n319_), .A2(G183gat), .A3(G190gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n333_), .A2(new_n334_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n331_), .A2(new_n332_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT25), .B(G183gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(G169gat), .B2(G176gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT78), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(G169gat), .B2(G176gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n341_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n340_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n328_), .B1(new_n337_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n351_));
  INV_X1    g150(.A(G211gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(G218gat), .ZN(new_n353_));
  INV_X1    g152(.A(G218gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(G211gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n351_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(G211gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(G218gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT88), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G197gat), .A2(G204gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(KEYINPUT21), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT21), .ZN(new_n365_));
  AND2_X1   g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(new_n366_), .B2(new_n361_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT87), .B(new_n365_), .C1(new_n366_), .C2(new_n361_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n360_), .A2(new_n364_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n364_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n359_), .A3(new_n356_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n350_), .A2(KEYINPUT92), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT92), .B1(new_n350_), .B2(new_n374_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT77), .B(G190gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(G183gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n318_), .B1(new_n337_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n359_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT88), .B1(new_n357_), .B2(new_n358_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n381_), .A2(new_n364_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n372_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n369_), .A2(new_n370_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n378_), .A2(KEYINPUT26), .ZN(new_n387_));
  NOR2_X1   g186(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n338_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n326_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n344_), .A2(new_n346_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n341_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n389_), .A2(new_n390_), .A3(new_n347_), .A4(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n380_), .A2(new_n386_), .A3(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n394_), .A2(KEYINPUT20), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n316_), .B1(new_n377_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G8gat), .B(G36gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT18), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n386_), .B1(new_n380_), .B2(new_n393_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT20), .B1(new_n350_), .B2(new_n374_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n316_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n396_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n400_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n350_), .A2(new_n374_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT92), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n350_), .A2(KEYINPUT92), .A3(new_n374_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(KEYINPUT20), .A3(new_n394_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n403_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n404_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n406_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n313_), .B1(new_n405_), .B2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n403_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n411_), .B2(new_n403_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n400_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(new_n413_), .A3(new_n406_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT27), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G78gat), .B(G106gat), .Z(new_n422_));
  INV_X1    g221(.A(KEYINPUT86), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT1), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n424_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT1), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(G155gat), .A3(G162gat), .ZN(new_n430_));
  OR2_X1    g229(.A1(G155gat), .A2(G162gat), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n427_), .A2(new_n428_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G141gat), .B(G148gat), .Z(new_n433_));
  INV_X1    g232(.A(KEYINPUT2), .ZN(new_n434_));
  INV_X1    g233(.A(G141gat), .ZN(new_n435_));
  INV_X1    g234(.A(G148gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n437_), .A2(new_n439_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n431_), .A2(new_n424_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n432_), .A2(new_n433_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT29), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n423_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT85), .B1(new_n424_), .B2(KEYINPUT1), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n433_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n442_), .A2(new_n443_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n446_), .A2(new_n374_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(KEYINPUT29), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n453_), .B1(new_n374_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n456_), .B2(KEYINPUT89), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n456_), .A2(KEYINPUT89), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n422_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n374_), .A2(new_n455_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(new_n461_), .B2(new_n453_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n456_), .A2(KEYINPUT89), .ZN(new_n463_));
  INV_X1    g262(.A(new_n422_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n454_), .A4(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT28), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n444_), .A2(new_n466_), .A3(new_n445_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n449_), .A2(new_n450_), .A3(new_n445_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT28), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G22gat), .B(G50gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(KEYINPUT90), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n459_), .A2(new_n465_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT90), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n467_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n471_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n475_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n482_), .B1(new_n459_), .B2(new_n465_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n421_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n486_));
  INV_X1    g285(.A(G127gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(G134gat), .ZN(new_n488_));
  INV_X1    g287(.A(G134gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(G127gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n486_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(G127gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(G134gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(KEYINPUT83), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G113gat), .B(G120gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n491_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n492_), .A2(new_n493_), .A3(KEYINPUT83), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT83), .B1(new_n492_), .B2(new_n493_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n451_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n496_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n444_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n503_), .A3(KEYINPUT4), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT93), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n501_), .A2(new_n503_), .A3(KEYINPUT93), .A4(KEYINPUT4), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n444_), .A2(new_n502_), .A3(KEYINPUT4), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G225gat), .A2(G233gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G1gat), .B(G29gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(G85gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT0), .B(G57gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n512_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n513_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n508_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n511_), .B1(new_n522_), .B2(new_n507_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n517_), .B1(new_n523_), .B2(new_n519_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n502_), .B(KEYINPUT31), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n380_), .A2(new_n393_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT30), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(G15gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G71gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n204_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n529_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n535_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT82), .B(G43gat), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n537_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n526_), .B(new_n528_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n526_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n541_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n539_), .A2(new_n535_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n530_), .A2(new_n536_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n537_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT84), .A3(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n545_), .A2(new_n551_), .A3(new_n527_), .ZN(new_n552_));
  AND4_X1   g351(.A1(new_n485_), .A2(new_n525_), .A3(new_n544_), .A4(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n415_), .A2(new_n484_), .A3(new_n420_), .A4(new_n525_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT97), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n521_), .A2(new_n524_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n556_), .A2(new_n477_), .A3(new_n483_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n415_), .A4(new_n420_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n406_), .A2(KEYINPUT32), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n417_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n412_), .A2(new_n413_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n560_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(new_n525_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT33), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n524_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n565_), .B1(new_n524_), .B2(new_n566_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n400_), .B1(new_n396_), .B2(new_n404_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT33), .B(new_n517_), .C1(new_n523_), .C2(new_n519_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT95), .B1(new_n501_), .B2(new_n503_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n511_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n501_), .A2(new_n503_), .A3(KEYINPUT95), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n517_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n512_), .B2(new_n510_), .ZN(new_n577_));
  AND4_X1   g376(.A1(new_n419_), .A2(new_n571_), .A3(new_n572_), .A4(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n564_), .B1(new_n570_), .B2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n555_), .B(new_n559_), .C1(new_n579_), .C2(new_n484_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n552_), .A2(new_n544_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n553_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n311_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT71), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n240_), .A2(new_n241_), .A3(new_n285_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n298_), .A2(new_n238_), .B1(new_n587_), .B2(new_n586_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(KEYINPUT71), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT73), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT37), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n599_), .B(KEYINPUT36), .Z(new_n606_));
  NAND3_X1  g405(.A1(new_n594_), .A2(new_n595_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n604_), .A3(KEYINPUT37), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n293_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(new_n253_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT74), .ZN(new_n617_));
  XOR2_X1   g416(.A(G127gat), .B(G155gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G183gat), .B(G211gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT17), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n617_), .A2(KEYINPUT75), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT75), .B1(new_n617_), .B2(new_n622_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT17), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n621_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n616_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n613_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n583_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n288_), .A3(new_n556_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT98), .B1(new_n311_), .B2(new_n630_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n582_), .A2(new_n609_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n280_), .A2(new_n638_), .A3(new_n629_), .A4(new_n310_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n636_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n288_), .B1(new_n640_), .B2(new_n556_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n635_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n634_), .B2(new_n633_), .ZN(G1324gat));
  NAND3_X1  g442(.A1(new_n632_), .A2(new_n289_), .A3(new_n421_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n636_), .A2(new_n421_), .A3(new_n637_), .A4(new_n639_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G8gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT99), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n649_), .A3(G8gat), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n647_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n648_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n644_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT40), .B(new_n644_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1325gat));
  INV_X1    g456(.A(new_n581_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n632_), .A2(new_n532_), .A3(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT100), .Z(new_n660_));
  NAND2_X1  g459(.A1(new_n640_), .A2(new_n658_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G15gat), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT41), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT41), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n660_), .A2(new_n663_), .A3(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n632_), .A2(new_n666_), .A3(new_n484_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n640_), .A2(new_n484_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G22gat), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n629_), .A2(new_n608_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n583_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT104), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n583_), .A2(new_n676_), .A3(new_n673_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(G29gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n556_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n555_), .A2(new_n559_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n569_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n578_), .A2(new_n682_), .A3(new_n567_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n563_), .A2(new_n525_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n484_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n581_), .B1(new_n681_), .B2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n581_), .A2(new_n556_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n485_), .ZN(new_n688_));
  AOI211_X1 g487(.A(KEYINPUT43), .B(new_n612_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n686_), .A2(new_n688_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n613_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT101), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n582_), .B2(new_n612_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n691_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n311_), .A2(new_n629_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(KEYINPUT44), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n556_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n698_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT102), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n701_), .A2(new_n705_), .A3(new_n702_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n700_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(new_n679_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n707_), .A2(KEYINPUT103), .A3(new_n679_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n680_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  INV_X1    g511(.A(new_n421_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(G36gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n675_), .A2(new_n677_), .A3(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT45), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n699_), .A2(new_n421_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n716_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n716_), .B(KEYINPUT46), .C1(new_n718_), .C2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1329gat));
  INV_X1    g523(.A(new_n699_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n726_));
  INV_X1    g525(.A(G43gat), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n581_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n678_), .A2(new_n658_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT47), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n729_), .A2(new_n734_), .A3(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1330gat));
  AOI21_X1  g535(.A(G50gat), .B1(new_n678_), .B2(new_n484_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n484_), .A2(G50gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n726_), .B2(new_n738_), .ZN(G1331gat));
  NOR3_X1   g538(.A1(new_n280_), .A2(new_n582_), .A3(new_n310_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n631_), .ZN(new_n741_));
  INV_X1    g540(.A(G57gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n556_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n310_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n625_), .A2(new_n628_), .A3(new_n744_), .ZN(new_n745_));
  NOR4_X1   g544(.A1(new_n280_), .A2(new_n582_), .A3(new_n609_), .A4(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(new_n556_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n742_), .B2(new_n747_), .ZN(G1332gat));
  INV_X1    g547(.A(G64gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n746_), .B2(new_n421_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT48), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n741_), .A2(new_n749_), .A3(new_n421_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1333gat));
  INV_X1    g552(.A(G71gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n746_), .B2(new_n658_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT105), .B(KEYINPUT49), .Z(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n741_), .A2(new_n754_), .A3(new_n658_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1334gat));
  INV_X1    g558(.A(G78gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n746_), .B2(new_n484_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT50), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n741_), .A2(new_n760_), .A3(new_n484_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1335gat));
  AND2_X1   g563(.A1(new_n740_), .A2(new_n673_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n556_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n696_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n694_), .A2(KEYINPUT101), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n691_), .A2(new_n695_), .A3(KEYINPUT106), .A4(new_n696_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT69), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n279_), .B(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n630_), .A3(new_n744_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT107), .B1(new_n772_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n778_), .B(new_n775_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n556_), .A2(new_n232_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n766_), .B1(new_n780_), .B2(new_n781_), .ZN(G1336gat));
  INV_X1    g581(.A(G92gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n765_), .A2(new_n783_), .A3(new_n421_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n777_), .A2(new_n779_), .A3(new_n713_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n783_), .ZN(G1337gat));
  AOI21_X1  g585(.A(new_n204_), .B1(new_n780_), .B2(new_n658_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n765_), .A2(new_n235_), .A3(new_n658_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT108), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  INV_X1    g590(.A(new_n789_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n777_), .A2(new_n779_), .A3(new_n581_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n791_), .B(new_n792_), .C1(new_n793_), .C2(new_n204_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(new_n794_), .ZN(G1338gat));
  OAI211_X1 g594(.A(new_n484_), .B(new_n776_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(G106gat), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  XOR2_X1   g598(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n797_), .A2(new_n798_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n484_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(G106gat), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n765_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  OR3_X1    g609(.A1(new_n804_), .A2(new_n808_), .A3(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(G1339gat));
  INV_X1    g612(.A(new_n745_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n279_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(KEYINPUT112), .A3(new_n279_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n612_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT54), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n817_), .A2(new_n821_), .A3(new_n612_), .A4(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n299_), .A2(new_n294_), .A3(new_n301_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n305_), .B1(new_n300_), .B2(new_n295_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n302_), .A2(new_n305_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n278_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT117), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n278_), .A2(new_n830_), .A3(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n310_), .A2(new_n277_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT12), .B1(new_n242_), .B2(new_n253_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n260_), .A2(new_n267_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT114), .B(new_n263_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n259_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n260_), .B(new_n267_), .C1(new_n839_), .C2(KEYINPUT12), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT114), .B1(new_n840_), .B2(new_n263_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n840_), .B2(new_n263_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n269_), .B2(new_n843_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n269_), .B2(new_n846_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n842_), .B(new_n845_), .C1(new_n847_), .C2(new_n849_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n850_), .A2(KEYINPUT56), .A3(new_n274_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT56), .B1(new_n850_), .B2(new_n274_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n834_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n832_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT116), .B(new_n834_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n609_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT57), .B1(new_n857_), .B2(KEYINPUT118), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n829_), .A2(new_n831_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n850_), .A2(new_n274_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n850_), .A2(KEYINPUT56), .A3(new_n274_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n833_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n859_), .B1(new_n864_), .B2(KEYINPUT116), .ZN(new_n865_));
  INV_X1    g664(.A(new_n856_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n608_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n277_), .B(new_n827_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n612_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n872_), .B2(new_n871_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n858_), .A2(new_n870_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n824_), .B1(new_n875_), .B2(new_n630_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n658_), .A2(new_n485_), .A3(new_n556_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G113gat), .B1(new_n878_), .B2(new_n310_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n853_), .A2(new_n854_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n856_), .A3(new_n859_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT118), .B1(new_n881_), .B2(new_n608_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n874_), .B1(new_n882_), .B2(new_n869_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n857_), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n630_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n823_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887_));
  INV_X1    g686(.A(new_n877_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(new_n878_), .B2(new_n887_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n886_), .A2(new_n888_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(KEYINPUT59), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n890_), .B1(new_n891_), .B2(new_n894_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n310_), .A2(G113gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n879_), .B1(new_n895_), .B2(new_n896_), .ZN(G1340gat));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n280_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n878_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n889_), .A2(new_n774_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n891_), .B2(new_n894_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n902_), .B2(new_n898_), .ZN(G1341gat));
  NOR3_X1   g702(.A1(new_n876_), .A2(new_n630_), .A3(new_n877_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT120), .B1(new_n904_), .B2(G127gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n886_), .A2(new_n629_), .A3(new_n888_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n487_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n630_), .A2(new_n487_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n895_), .B2(new_n910_), .ZN(G1342gat));
  AOI21_X1  g710(.A(G134gat), .B1(new_n878_), .B2(new_n609_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n613_), .A2(G134gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT121), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n895_), .B2(new_n914_), .ZN(G1343gat));
  NAND3_X1  g714(.A1(new_n713_), .A2(new_n484_), .A3(new_n556_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n876_), .A2(new_n658_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n310_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT122), .B(G141gat), .Z(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1344gat));
  NAND2_X1  g719(.A1(new_n917_), .A2(new_n774_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g721(.A1(new_n917_), .A2(new_n629_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT61), .B(G155gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1346gat));
  AOI21_X1  g724(.A(G162gat), .B1(new_n917_), .B2(new_n609_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n613_), .A2(G162gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT123), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n917_), .B2(new_n928_), .ZN(G1347gat));
  INV_X1    g728(.A(G169gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n687_), .A2(new_n805_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n886_), .A2(new_n421_), .A3(new_n310_), .A4(new_n934_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n930_), .B(new_n932_), .C1(new_n935_), .C2(KEYINPUT22), .ZN(new_n936_));
  NOR4_X1   g735(.A1(new_n876_), .A2(new_n713_), .A3(new_n744_), .A4(new_n933_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT22), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n931_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(G169gat), .B1(new_n935_), .B2(new_n932_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n936_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(G1348gat));
  NAND4_X1  g741(.A1(new_n886_), .A2(new_n421_), .A3(new_n774_), .A4(new_n934_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g743(.A1(new_n886_), .A2(new_n629_), .A3(new_n421_), .A4(new_n934_), .ZN(new_n945_));
  MUX2_X1   g744(.A(new_n338_), .B(G183gat), .S(new_n945_), .Z(G1350gat));
  NAND2_X1  g745(.A1(new_n886_), .A2(new_n421_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n933_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n948_), .A2(new_n609_), .A3(new_n339_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n947_), .A2(new_n612_), .A3(new_n933_), .ZN(new_n950_));
  INV_X1    g749(.A(G190gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n949_), .B1(new_n950_), .B2(new_n951_), .ZN(G1351gat));
  AND4_X1   g751(.A1(new_n421_), .A2(new_n886_), .A3(new_n581_), .A4(new_n557_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(new_n310_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(KEYINPUT125), .B(G197gat), .ZN(new_n955_));
  INV_X1    g754(.A(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n956_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n953_), .A2(new_n310_), .A3(new_n955_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1352gat));
  NAND2_X1  g758(.A1(new_n953_), .A2(new_n774_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(G204gat), .ZN(new_n961_));
  INV_X1    g760(.A(G204gat), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n953_), .A2(new_n962_), .A3(new_n774_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n963_), .ZN(G1353gat));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n629_), .B1(new_n965_), .B2(new_n352_), .ZN(new_n966_));
  XOR2_X1   g765(.A(new_n966_), .B(KEYINPUT126), .Z(new_n967_));
  NAND3_X1  g766(.A1(new_n965_), .A2(new_n352_), .A3(KEYINPUT127), .ZN(new_n968_));
  AND3_X1   g767(.A1(new_n953_), .A2(new_n967_), .A3(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n970_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n971_));
  AOI22_X1  g770(.A1(new_n953_), .A2(new_n967_), .B1(new_n971_), .B2(new_n968_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n969_), .A2(new_n972_), .ZN(G1354gat));
  NAND3_X1  g772(.A1(new_n953_), .A2(new_n354_), .A3(new_n609_), .ZN(new_n974_));
  AND2_X1   g773(.A1(new_n953_), .A2(new_n613_), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n974_), .B1(new_n975_), .B2(new_n354_), .ZN(G1355gat));
endmodule


