//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n205_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G229gat), .A2(G233gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n204_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n212_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n212_), .B2(new_n205_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n216_), .B1(new_n220_), .B2(new_n215_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G113gat), .B(G141gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G169gat), .B(G197gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n222_), .B(new_n223_), .Z(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT76), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n225_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT6), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT65), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT6), .ZN(new_n235_));
  AND2_X1   g034(.A1(G99gat), .A2(G106gat), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n233_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n236_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n240_));
  INV_X1    g039(.A(G106gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT9), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT64), .B(G85gat), .ZN(new_n247_));
  INV_X1    g046(.A(G92gat), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(KEYINPUT9), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n243_), .B(new_n246_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n239_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT7), .ZN(new_n253_));
  INV_X1    g052(.A(G99gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n241_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G99gat), .A2(G106gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n234_), .A2(KEYINPUT6), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n232_), .A2(KEYINPUT65), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n233_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n257_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n244_), .A2(new_n245_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n263_), .A2(KEYINPUT8), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT8), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n255_), .A2(new_n256_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n267_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n264_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n266_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n252_), .B1(new_n265_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT8), .B1(new_n263_), .B2(new_n264_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n268_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n251_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT66), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT11), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G71gat), .B(G78gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n279_), .A2(new_n280_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT11), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n279_), .A2(new_n280_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n282_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n281_), .A2(KEYINPUT11), .A3(new_n283_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT12), .B1(new_n278_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n290_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n273_), .A2(new_n277_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(KEYINPUT12), .A3(new_n271_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G230gat), .A2(G233gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n298_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n293_), .B1(new_n273_), .B2(new_n277_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n294_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  AOI211_X1 g102(.A(new_n272_), .B(new_n251_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n274_), .A2(new_n275_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT66), .B1(new_n305_), .B2(new_n252_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n291_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n307_), .A2(KEYINPUT68), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n300_), .B1(new_n303_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G120gat), .B(G148gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT5), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G176gat), .B(G204gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n299_), .A2(new_n309_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n299_), .B2(new_n309_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT13), .ZN(new_n317_));
  OR3_X1    g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n317_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(KEYINPUT69), .A3(new_n319_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n231_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT84), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G227gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(G15gat), .ZN(new_n328_));
  INV_X1    g127(.A(G71gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(new_n254_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G169gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G183gat), .A3(G190gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT81), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT79), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(G183gat), .A3(G190gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT23), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT80), .A4(KEYINPUT23), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n337_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(KEYINPUT77), .B(G190gat), .Z(new_n347_));
  INV_X1    g146(.A(G183gat), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n334_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT25), .B(G183gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n351_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT23), .B1(new_n339_), .B2(new_n341_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n335_), .B1(G183gat), .B2(G190gat), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT24), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(G169gat), .B2(G176gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT78), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(G169gat), .B2(G176gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n364_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n359_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n355_), .A2(new_n358_), .A3(new_n365_), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n350_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n350_), .A2(KEYINPUT30), .A3(new_n368_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n332_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n332_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT82), .B(G43gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n326_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(KEYINPUT84), .A3(new_n377_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G113gat), .B(G120gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G134gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G127gat), .ZN(new_n386_));
  INV_X1    g185(.A(G127gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G134gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n388_), .A3(KEYINPUT83), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT83), .B1(new_n386_), .B2(new_n388_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n384_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n386_), .A2(new_n388_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n389_), .A3(new_n383_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT31), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n380_), .A2(new_n382_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT1), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT1), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(G155gat), .A3(G162gat), .ZN(new_n408_));
  OR2_X1    g207(.A1(G155gat), .A2(G162gat), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n405_), .A2(new_n406_), .A3(new_n408_), .A4(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G141gat), .B(G148gat), .Z(new_n411_));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412_));
  INV_X1    g211(.A(G141gat), .ZN(new_n413_));
  INV_X1    g212(.A(G148gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G141gat), .A2(G148gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT2), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n415_), .A2(new_n418_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n409_), .A2(new_n402_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n410_), .A2(new_n411_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n397_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n406_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT85), .B1(new_n402_), .B2(KEYINPUT1), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n411_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n421_), .A2(new_n422_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(new_n396_), .A3(new_n392_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n401_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n424_), .A2(new_n430_), .A3(KEYINPUT4), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n424_), .A2(new_n430_), .A3(KEYINPUT93), .A4(KEYINPUT4), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n430_), .A2(KEYINPUT4), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n431_), .B1(new_n438_), .B2(new_n401_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G85gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT0), .B(G57gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n436_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n400_), .B1(new_n446_), .B2(new_n435_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n443_), .B1(new_n447_), .B2(new_n431_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n398_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n326_), .B(new_n450_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G197gat), .B(G204gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT21), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G218gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(G211gat), .ZN(new_n456_));
  INV_X1    g255(.A(G211gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G218gat), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n456_), .A2(new_n458_), .A3(KEYINPUT88), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT88), .B1(new_n456_), .B2(new_n458_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n454_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n452_), .A2(new_n453_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  OAI221_X1 g265(.A(new_n454_), .B1(new_n459_), .B2(new_n460_), .C1(new_n464_), .C2(new_n462_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n429_), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT29), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n423_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G228gat), .A2(G233gat), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n469_), .A2(new_n470_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n466_), .B(new_n467_), .C1(new_n472_), .C2(new_n423_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n477_));
  INV_X1    g276(.A(new_n474_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n475_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G78gat), .B(G106gat), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G22gat), .B(G50gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT28), .B1(new_n429_), .B2(KEYINPUT29), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT28), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n423_), .A2(new_n486_), .A3(new_n472_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n484_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(new_n487_), .A3(new_n484_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT90), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n482_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n475_), .B(new_n493_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n483_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496_));
  INV_X1    g295(.A(new_n490_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n488_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(new_n483_), .B2(new_n494_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n399_), .A2(new_n449_), .A3(new_n451_), .A4(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT96), .B(KEYINPUT27), .ZN(new_n504_));
  OAI22_X1  g303(.A1(new_n356_), .A2(new_n357_), .B1(G183gat), .B2(G190gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n334_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT26), .B(G190gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n351_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n361_), .A2(new_n359_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n365_), .A3(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n506_), .B1(new_n346_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n469_), .A2(KEYINPUT92), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n344_), .A2(new_n345_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n337_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n510_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n516_), .A2(new_n517_), .B1(new_n334_), .B2(new_n505_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n513_), .B1(new_n518_), .B2(new_n468_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n350_), .A2(new_n468_), .A3(new_n368_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n512_), .A2(new_n519_), .A3(KEYINPUT20), .A4(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G226gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT20), .B1(new_n469_), .B2(new_n511_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n468_), .B1(new_n350_), .B2(new_n368_), .ZN(new_n528_));
  OR3_X1    g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n525_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G8gat), .B(G36gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT18), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G64gat), .B(G92gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  AND3_X1   g332(.A1(new_n526_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n504_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n525_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n521_), .B2(new_n525_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n533_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n526_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(KEYINPUT27), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n503_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n483_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n500_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n449_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT97), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n445_), .A2(new_n448_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n549_), .A2(new_n495_), .A3(new_n500_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT97), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(new_n536_), .A4(new_n542_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n533_), .A2(KEYINPUT32), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n526_), .A2(new_n529_), .A3(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n538_), .A2(KEYINPUT32), .A3(new_n533_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n549_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT33), .B(new_n443_), .C1(new_n447_), .C2(new_n431_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n424_), .A2(new_n430_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n400_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(new_n560_), .B2(new_n559_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n562_), .B(new_n444_), .C1(new_n438_), .C2(new_n401_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n564_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT33), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n566_), .B(new_n567_), .C1(new_n439_), .C2(new_n444_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n566_), .B1(new_n448_), .B2(new_n567_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n557_), .B1(new_n565_), .B2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n548_), .B(new_n552_), .C1(new_n572_), .C2(new_n501_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n399_), .A2(new_n451_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n544_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n212_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n293_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT74), .ZN(new_n579_));
  XOR2_X1   g378(.A(G127gat), .B(G155gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G183gat), .B(G211gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT17), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT75), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n578_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n304_), .A2(new_n306_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n204_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n218_), .A2(new_n271_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT34), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT71), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n601_), .B2(new_n605_), .ZN(new_n609_));
  AOI211_X1 g408(.A(KEYINPUT71), .B(new_n604_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n610_));
  OAI221_X1 g409(.A(new_n597_), .B1(new_n601_), .B2(new_n607_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n601_), .A2(new_n607_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n595_), .B(KEYINPUT36), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT73), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n611_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  OAI221_X1 g419(.A(new_n611_), .B1(new_n618_), .B2(new_n617_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR4_X1   g422(.A1(new_n325_), .A2(new_n575_), .A3(new_n592_), .A4(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n207_), .A3(new_n549_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT38), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT98), .B1(new_n325_), .B2(new_n592_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n324_), .A2(new_n628_), .A3(new_n591_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n616_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n575_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n627_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n449_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n633_), .ZN(G1324gat));
  NAND3_X1  g433(.A1(new_n624_), .A2(new_n208_), .A3(new_n543_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n543_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G8gat), .B1(new_n632_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT99), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n640_), .B(G8gat), .C1(new_n632_), .C2(new_n636_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n639_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n635_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT40), .B(new_n635_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n632_), .B2(new_n574_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT41), .Z(new_n650_));
  INV_X1    g449(.A(G15gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n574_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n624_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT100), .Z(new_n654_));
  NAND2_X1  g453(.A1(new_n650_), .A2(new_n654_), .ZN(G1326gat));
  OAI21_X1  g454(.A(G22gat), .B1(new_n632_), .B2(new_n502_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT42), .ZN(new_n657_));
  INV_X1    g456(.A(G22gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n624_), .A2(new_n658_), .A3(new_n501_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1327gat));
  NOR2_X1   g459(.A1(new_n325_), .A2(new_n575_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n591_), .A2(new_n616_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(KEYINPUT104), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(KEYINPUT104), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OR3_X1    g465(.A1(new_n666_), .A2(G29gat), .A3(new_n449_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n325_), .A2(new_n591_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n548_), .A2(new_n552_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n565_), .A2(new_n571_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n501_), .B1(new_n670_), .B2(new_n556_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n574_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n544_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n623_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT101), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n674_), .A2(new_n679_), .A3(new_n675_), .A4(new_n623_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT43), .B1(new_n575_), .B2(new_n622_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT44), .B(new_n668_), .C1(new_n678_), .C2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n668_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n680_), .A2(new_n681_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n677_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n686_), .A2(KEYINPUT102), .A3(KEYINPUT44), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n668_), .B1(new_n678_), .B2(new_n682_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n549_), .B(new_n683_), .C1(new_n687_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G29gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n667_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(new_n683_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT102), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n689_), .A2(new_n688_), .A3(new_n690_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n698_), .B1(new_n702_), .B2(new_n543_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n636_), .A2(G36gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n664_), .A2(new_n665_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT45), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n664_), .A2(new_n707_), .A3(new_n665_), .A4(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n697_), .B1(new_n703_), .B2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n543_), .B(new_n683_), .C1(new_n687_), .C2(new_n691_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G36gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(KEYINPUT46), .A3(new_n709_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1329gat));
  INV_X1    g514(.A(G43gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n574_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n702_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n666_), .B2(new_n574_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT47), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n718_), .A2(new_n722_), .A3(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1330gat));
  INV_X1    g523(.A(new_n666_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G50gat), .B1(new_n725_), .B2(new_n501_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n501_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n702_), .B2(new_n727_), .ZN(G1331gat));
  NAND2_X1  g527(.A1(new_n322_), .A2(new_n323_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n575_), .A2(new_n729_), .A3(new_n230_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n730_), .A2(new_n591_), .A3(new_n622_), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n549_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n591_), .A3(new_n616_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n449_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1332gat));
  OAI21_X1  g535(.A(G64gat), .B1(new_n734_), .B2(new_n636_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT48), .ZN(new_n738_));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n731_), .A2(new_n739_), .A3(new_n543_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1333gat));
  NAND3_X1  g540(.A1(new_n731_), .A2(new_n329_), .A3(new_n652_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n734_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n329_), .B1(new_n743_), .B2(new_n652_), .ZN(new_n744_));
  XOR2_X1   g543(.A(KEYINPUT105), .B(KEYINPUT49), .Z(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n744_), .A2(new_n745_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n742_), .B1(new_n747_), .B2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n734_), .B2(new_n502_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n731_), .A2(new_n752_), .A3(new_n501_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1335gat));
  AND2_X1   g553(.A1(new_n730_), .A2(new_n662_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n549_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n677_), .A2(new_n681_), .A3(new_n758_), .A4(new_n680_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n729_), .A2(new_n591_), .A3(new_n230_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n758_), .B1(new_n685_), .B2(new_n677_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT106), .B1(new_n678_), .B2(new_n682_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n764_), .A2(KEYINPUT107), .A3(new_n759_), .A4(new_n760_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n449_), .A2(new_n247_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n756_), .B1(new_n766_), .B2(new_n767_), .ZN(G1336gat));
  NAND3_X1  g567(.A1(new_n755_), .A2(new_n248_), .A3(new_n543_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n766_), .A2(new_n543_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n248_), .ZN(G1337gat));
  NAND3_X1  g570(.A1(new_n763_), .A2(new_n652_), .A3(new_n765_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G99gat), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n652_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n755_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT51), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n773_), .A2(new_n779_), .A3(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1338gat));
  OAI211_X1 g580(.A(new_n501_), .B(new_n760_), .C1(new_n678_), .C2(new_n682_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783_));
  XOR2_X1   g582(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n782_), .A2(new_n783_), .A3(G106gat), .A4(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n755_), .A2(new_n241_), .A3(new_n501_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n785_), .A2(new_n783_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n784_), .A2(KEYINPUT110), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n789_), .B(new_n790_), .C1(new_n782_), .C2(G106gat), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n788_), .A2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1339gat));
  NOR2_X1   g593(.A1(new_n574_), .A2(new_n501_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n543_), .A2(new_n449_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n294_), .B(new_n295_), .C1(new_n301_), .C2(KEYINPUT12), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n300_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n800_), .B(new_n300_), .C1(new_n292_), .C2(new_n296_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n798_), .B2(new_n300_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n297_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n298_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT12), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n293_), .A2(new_n276_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n598_), .B2(new_n293_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n307_), .A2(new_n806_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(KEYINPUT55), .A4(new_n298_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n805_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n313_), .B1(new_n804_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n315_), .B1(new_n814_), .B2(KEYINPUT56), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n313_), .C1(new_n804_), .C2(new_n813_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n224_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n220_), .B2(new_n214_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n226_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n815_), .A2(KEYINPUT58), .A3(new_n817_), .A4(new_n820_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n623_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n814_), .A2(KEYINPUT56), .ZN(new_n827_));
  INV_X1    g626(.A(new_n315_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n230_), .A3(new_n828_), .A4(new_n817_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n815_), .A2(KEYINPUT116), .A3(new_n230_), .A4(new_n817_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n820_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT117), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n835_), .B(new_n820_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n831_), .A2(new_n832_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n616_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n826_), .B1(new_n842_), .B2(KEYINPUT57), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n840_), .A2(new_n841_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n591_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n591_), .A2(new_n231_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n320_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(KEYINPUT112), .A3(new_n591_), .A4(new_n231_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n622_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT54), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n849_), .A2(new_n854_), .A3(new_n851_), .A4(new_n622_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n795_), .B(new_n796_), .C1(new_n846_), .C2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G113gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n230_), .ZN(new_n860_));
  OR2_X1    g659(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n861_));
  NAND2_X1  g660(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n796_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n837_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n630_), .B1(new_n865_), .B2(new_n832_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT57), .B1(new_n866_), .B2(KEYINPUT118), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n845_), .A2(new_n867_), .A3(new_n825_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n592_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n856_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n864_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n871_), .A2(KEYINPUT119), .A3(KEYINPUT59), .A4(new_n795_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n231_), .B1(new_n863_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n860_), .B1(new_n873_), .B2(new_n859_), .ZN(G1340gat));
  INV_X1    g673(.A(G120gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n729_), .B2(KEYINPUT60), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n858_), .B(new_n876_), .C1(KEYINPUT60), .C2(new_n875_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n729_), .B1(new_n863_), .B2(new_n872_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n875_), .ZN(G1341gat));
  AOI21_X1  g678(.A(new_n856_), .B1(new_n868_), .B2(new_n592_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n795_), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n880_), .A2(new_n592_), .A3(new_n881_), .A4(new_n864_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT120), .B1(new_n882_), .B2(G127gat), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n884_), .B(new_n387_), .C1(new_n857_), .C2(new_n592_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n591_), .A2(G127gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n863_), .B2(new_n872_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1342gat));
  AOI21_X1  g688(.A(G134gat), .B1(new_n858_), .B2(new_n630_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n863_), .A2(new_n872_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n623_), .A2(G134gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT121), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n891_), .B2(new_n893_), .ZN(G1343gat));
  NOR2_X1   g693(.A1(new_n652_), .A2(new_n502_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n871_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n230_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT122), .B(G141gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n896_), .A2(new_n230_), .A3(new_n898_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1344gat));
  INV_X1    g701(.A(new_n729_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n896_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G148gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n896_), .A2(new_n414_), .A3(new_n903_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1345gat));
  NAND2_X1  g706(.A1(new_n896_), .A2(new_n591_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G155gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n909_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n896_), .A2(new_n591_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n896_), .B2(new_n630_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n623_), .A2(G162gat), .ZN(new_n915_));
  XOR2_X1   g714(.A(new_n915_), .B(KEYINPUT123), .Z(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n896_), .B2(new_n916_), .ZN(G1347gat));
  NOR4_X1   g716(.A1(new_n880_), .A2(new_n231_), .A3(new_n636_), .A4(new_n503_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT22), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n920_), .A2(G169gat), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n924_));
  INV_X1    g723(.A(G169gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n918_), .B2(new_n921_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n923_), .B1(new_n924_), .B2(new_n926_), .ZN(G1348gat));
  NOR2_X1   g726(.A1(new_n880_), .A2(new_n636_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n503_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n928_), .A2(new_n903_), .A3(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g730(.A1(new_n928_), .A2(new_n591_), .A3(new_n929_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n351_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n933_), .B1(new_n348_), .B2(new_n932_), .ZN(G1350gat));
  NAND2_X1  g733(.A1(new_n928_), .A2(new_n929_), .ZN(new_n935_));
  OAI21_X1  g734(.A(G190gat), .B1(new_n935_), .B2(new_n622_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n630_), .A2(new_n507_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n935_), .B2(new_n937_), .ZN(G1351gat));
  NAND2_X1  g737(.A1(new_n895_), .A2(new_n449_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n880_), .A2(new_n636_), .A3(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n230_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT125), .B(G197gat), .ZN(new_n942_));
  XOR2_X1   g741(.A(new_n941_), .B(new_n942_), .Z(G1352gat));
  NAND2_X1  g742(.A1(new_n940_), .A2(new_n903_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g744(.A(new_n592_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT126), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n940_), .A2(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n949_), .A2(KEYINPUT127), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(KEYINPUT127), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n948_), .A2(new_n950_), .A3(new_n951_), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n940_), .A2(KEYINPUT127), .A3(new_n947_), .A4(new_n949_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1354gat));
  NAND3_X1  g753(.A1(new_n940_), .A2(new_n455_), .A3(new_n630_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n940_), .A2(new_n623_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n455_), .ZN(G1355gat));
endmodule


