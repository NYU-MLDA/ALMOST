//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n203_));
  OAI211_X1 g002(.A(G85gat), .B(G92gat), .C1(new_n203_), .C2(KEYINPUT9), .ZN(new_n204_));
  OAI211_X1 g003(.A(new_n203_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT65), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(KEYINPUT65), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT10), .B(G99gat), .Z(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n207_), .A2(new_n209_), .A3(new_n210_), .A4(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n209_), .A2(KEYINPUT66), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT7), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n209_), .A2(KEYINPUT66), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G85gat), .B(G92gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n215_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  AOI211_X1 g022(.A(KEYINPUT8), .B(new_n221_), .C1(new_n218_), .C2(new_n209_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n214_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G57gat), .B(G64gat), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(KEYINPUT11), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(KEYINPUT11), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G78gat), .Z(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n228_), .A2(new_n229_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n225_), .A2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n214_), .B(new_n232_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(KEYINPUT12), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT12), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n225_), .A2(new_n237_), .A3(new_n233_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G230gat), .A2(G233gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n234_), .A2(new_n235_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n240_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G120gat), .B(G148gat), .Z(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G176gat), .B(G204gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n241_), .A2(new_n244_), .A3(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(KEYINPUT13), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT13), .B1(new_n251_), .B2(new_n253_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n202_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT68), .A3(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G29gat), .B(G36gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G43gat), .B(G50gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT15), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT35), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G232gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT34), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n225_), .A2(new_n264_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n265_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n214_), .B(new_n263_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n269_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n271_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G190gat), .B(G218gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G134gat), .B(G162gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NOR4_X1   g077(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT36), .A4(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(KEYINPUT36), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n275_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(new_n273_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT37), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT69), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT69), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(KEYINPUT69), .B(new_n285_), .C1(new_n279_), .C2(new_n283_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT71), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n232_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G8gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G15gat), .ZN(new_n297_));
  INV_X1    g096(.A(G22gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G15gat), .A2(G22gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G1gat), .A2(G8gat), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n299_), .A2(new_n300_), .B1(KEYINPUT14), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n296_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n293_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT17), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G155gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT16), .ZN(new_n307_));
  XOR2_X1   g106(.A(G183gat), .B(G211gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n304_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(KEYINPUT17), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n304_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n290_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n260_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G113gat), .B(G141gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT73), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G169gat), .B(G197gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n303_), .B(new_n263_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G229gat), .A2(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n303_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n264_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n303_), .A2(new_n263_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n324_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n322_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  AOI211_X1 g132(.A(KEYINPUT74), .B(new_n321_), .C1(new_n326_), .C2(new_n330_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT75), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n333_), .A2(new_n334_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G211gat), .B(G218gat), .Z(new_n341_));
  NOR2_X1   g140(.A1(G197gat), .A2(G204gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n341_), .A2(KEYINPUT21), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(KEYINPUT21), .A3(new_n344_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT21), .ZN(new_n347_));
  AND2_X1   g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(new_n342_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n345_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353_));
  INV_X1    g152(.A(G155gat), .ZN(new_n354_));
  INV_X1    g153(.A(G162gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G141gat), .A2(G148gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT2), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n358_), .A2(KEYINPUT1), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G155gat), .A3(G162gat), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n356_), .A2(new_n369_), .A3(new_n371_), .A4(new_n357_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G141gat), .B(G148gat), .Z(new_n373_));
  AOI22_X1  g172(.A1(new_n359_), .A2(new_n368_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n352_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n352_), .B2(KEYINPUT85), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  OAI221_X1 g178(.A(new_n352_), .B1(KEYINPUT85), .B2(new_n377_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT87), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT87), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n379_), .A2(new_n380_), .A3(new_n385_), .A4(new_n382_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n382_), .B(KEYINPUT86), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n381_), .A2(KEYINPUT88), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G22gat), .B(G50gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n359_), .A2(new_n368_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n372_), .A2(new_n373_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT28), .B1(new_n394_), .B2(KEYINPUT29), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n394_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n391_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n397_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n395_), .A3(new_n390_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n387_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n398_), .B(new_n400_), .C1(new_n402_), .C2(KEYINPUT88), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n381_), .A2(new_n387_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(new_n402_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n398_), .A2(new_n400_), .ZN(new_n406_));
  OAI22_X1  g205(.A1(new_n389_), .A2(new_n403_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G127gat), .B(G134gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G113gat), .B(G120gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G134gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G127gat), .ZN(new_n414_));
  INV_X1    g213(.A(G127gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G134gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G120gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G113gat), .ZN(new_n419_));
  INV_X1    g218(.A(G113gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G120gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n422_), .A3(KEYINPUT81), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n410_), .A2(new_n411_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n412_), .B(new_n423_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT76), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G169gat), .A2(G176gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT24), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G183gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT25), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT25), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G183gat), .ZN(new_n437_));
  INV_X1    g236(.A(G190gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT26), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT26), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G190gat), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n435_), .A2(new_n437_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(G169gat), .ZN(new_n443_));
  INV_X1    g242(.A(G176gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n445_), .A2(KEYINPUT76), .A3(KEYINPUT24), .A4(new_n430_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n433_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT77), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT77), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n433_), .A2(new_n442_), .A3(new_n449_), .A4(new_n446_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT24), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n432_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n448_), .A2(new_n450_), .A3(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT79), .B(G176gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G169gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n443_), .A2(KEYINPUT78), .A3(KEYINPUT22), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n458_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n434_), .A2(new_n438_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n452_), .A2(new_n463_), .A3(new_n455_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n430_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n457_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G227gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(new_n297_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G99gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G71gat), .ZN(new_n471_));
  INV_X1    g270(.A(G71gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G99gat), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n471_), .A2(new_n473_), .A3(G43gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(G43gat), .B1(new_n471_), .B2(new_n473_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT30), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n477_));
  INV_X1    g276(.A(G43gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n472_), .A2(G99gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n470_), .A2(G71gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n471_), .A2(new_n473_), .A3(G43gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n477_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n469_), .B1(new_n476_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT30), .B1(new_n474_), .B2(new_n475_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n468_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n428_), .B1(new_n466_), .B2(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n485_), .A2(new_n468_), .A3(new_n486_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n468_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n465_), .ZN(new_n493_));
  AND3_X1   g292(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(new_n451_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n454_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n447_), .B2(KEYINPUT77), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n493_), .B1(new_n497_), .B2(new_n450_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n492_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT83), .B1(new_n489_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT31), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT82), .B1(new_n492_), .B2(new_n498_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT83), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n466_), .A2(new_n488_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n500_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n501_), .B1(new_n500_), .B2(new_n505_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n427_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n489_), .A2(new_n499_), .A3(KEYINPUT83), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n503_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT31), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n427_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n500_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n417_), .A2(new_n422_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n410_), .A2(new_n411_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n392_), .B(new_n393_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n427_), .B2(new_n374_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT4), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G225gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT92), .Z(new_n521_));
  AND2_X1   g320(.A1(new_n412_), .A2(new_n423_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT80), .B1(new_n417_), .B2(new_n422_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n410_), .A2(new_n411_), .A3(new_n424_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n522_), .A2(new_n394_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT4), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n519_), .A2(new_n521_), .A3(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G1gat), .B(G29gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G85gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT0), .B(G57gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n521_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n518_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n533_), .B1(new_n529_), .B2(new_n535_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n508_), .A2(new_n514_), .A3(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n345_), .A2(new_n351_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT22), .B(G169gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n458_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(new_n464_), .A3(new_n430_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n445_), .A2(KEYINPUT24), .A3(new_n430_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n442_), .A2(new_n495_), .A3(new_n545_), .A4(new_n454_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT20), .B(new_n547_), .C1(new_n498_), .C2(new_n541_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G226gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT19), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT94), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n546_), .A2(KEYINPUT90), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT25), .B(G183gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(G190gat), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n453_), .B1(G169gat), .B2(G176gat), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n557_), .A2(new_n558_), .B1(new_n559_), .B2(new_n445_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n556_), .B1(new_n560_), .B2(new_n456_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n544_), .B1(new_n555_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n352_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n457_), .A2(new_n465_), .A3(new_n541_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n550_), .B(KEYINPUT89), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(KEYINPUT20), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT95), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n562_), .B2(new_n352_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n565_), .A4(new_n564_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n552_), .A2(new_n554_), .B1(new_n567_), .B2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G8gat), .B(G36gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT18), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G64gat), .B(G92gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT96), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT97), .B1(new_n572_), .B2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n566_), .A2(KEYINPUT95), .ZN(new_n580_));
  INV_X1    g379(.A(new_n571_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n548_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n553_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n583_));
  OAI22_X1  g382(.A1(new_n580_), .A2(new_n581_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT97), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n577_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n541_), .B(new_n544_), .C1(new_n555_), .C2(new_n561_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT91), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n544_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n546_), .A2(KEYINPUT90), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n560_), .A2(new_n556_), .A3(new_n456_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT91), .A3(new_n541_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n589_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n550_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n568_), .B1(new_n466_), .B2(new_n352_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n565_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n564_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT20), .B1(new_n593_), .B2(new_n541_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(new_n576_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT27), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n579_), .A2(new_n586_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT27), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n598_), .A2(new_n576_), .A3(new_n602_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n576_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  AND4_X1   g409(.A1(new_n408_), .A2(new_n540_), .A3(new_n606_), .A4(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n508_), .A2(new_n514_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n598_), .A2(new_n602_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n576_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT27), .B1(new_n616_), .B2(new_n603_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n407_), .A2(new_n539_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n606_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n529_), .A2(new_n535_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n533_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n536_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n576_), .A2(KEYINPUT32), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n598_), .A2(new_n625_), .A3(new_n602_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n624_), .B(new_n626_), .C1(new_n572_), .C2(new_n625_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n533_), .B1(new_n518_), .B2(new_n534_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n519_), .A2(new_n528_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n629_), .B2(new_n534_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(KEYINPUT33), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n630_), .B1(new_n538_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n535_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n527_), .B1(new_n526_), .B2(new_n517_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT4), .B1(new_n512_), .B2(new_n394_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n635_), .B1(new_n638_), .B2(new_n521_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n632_), .B1(new_n639_), .B2(new_n533_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n616_), .A2(new_n634_), .A3(new_n640_), .A4(new_n603_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n627_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n408_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n613_), .B1(new_n620_), .B2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n611_), .B1(new_n644_), .B2(KEYINPUT98), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n606_), .A2(new_n619_), .B1(new_n642_), .B2(new_n408_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(new_n613_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n340_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n260_), .A2(KEYINPUT72), .A3(new_n314_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n317_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT99), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT99), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n539_), .A2(G1gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT38), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n652_), .A2(KEYINPUT38), .A3(new_n653_), .A4(new_n654_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n284_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT100), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(KEYINPUT100), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n260_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n663_), .A2(new_n335_), .A3(new_n313_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n624_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G1gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n658_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1324gat));
  NAND2_X1  g468(.A1(new_n584_), .A2(new_n577_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n604_), .B1(new_n670_), .B2(KEYINPUT97), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n617_), .B1(new_n671_), .B2(new_n586_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(G8gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n652_), .A2(new_n653_), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n675_));
  INV_X1    g474(.A(new_n672_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n664_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G8gat), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(KEYINPUT39), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(KEYINPUT39), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n674_), .B(new_n675_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n678_), .B(KEYINPUT39), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n675_), .B1(new_n683_), .B2(new_n674_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1325gat));
  INV_X1    g484(.A(new_n651_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n297_), .A3(new_n613_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n662_), .A2(new_n613_), .A3(new_n664_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n688_), .B2(G15gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(G1326gat));
  NAND3_X1  g490(.A1(new_n686_), .A2(new_n298_), .A3(new_n407_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n662_), .A2(new_n407_), .A3(new_n664_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G22gat), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT42), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(KEYINPUT42), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(G1327gat));
  INV_X1    g496(.A(new_n284_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n312_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n260_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(new_n649_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G29gat), .B1(new_n701_), .B2(new_n624_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n704_));
  INV_X1    g503(.A(new_n290_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n706_));
  XOR2_X1   g505(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n611_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n610_), .A2(new_n407_), .A3(new_n539_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n586_), .B2(new_n671_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n407_), .B1(new_n627_), .B2(new_n641_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT98), .B(new_n612_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n648_), .A2(new_n709_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n290_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n707_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(KEYINPUT104), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n714_), .A2(new_n718_), .A3(new_n290_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n714_), .A2(KEYINPUT105), .A3(new_n718_), .A4(new_n290_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n708_), .A2(new_n717_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n663_), .A2(new_n335_), .A3(new_n312_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n703_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT104), .B1(new_n715_), .B2(new_n716_), .ZN(new_n727_));
  AOI211_X1 g526(.A(new_n704_), .B(new_n707_), .C1(new_n714_), .C2(new_n290_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT105), .B1(new_n706_), .B2(new_n718_), .ZN(new_n729_));
  AND4_X1   g528(.A1(KEYINPUT105), .A2(new_n714_), .A3(new_n718_), .A4(new_n290_), .ZN(new_n730_));
  OAI22_X1  g529(.A1(new_n727_), .A2(new_n728_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(KEYINPUT44), .A3(new_n724_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n726_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n624_), .A2(G29gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n702_), .B1(new_n733_), .B2(new_n734_), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n726_), .A2(new_n732_), .A3(new_n676_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G36gat), .ZN(new_n737_));
  INV_X1    g536(.A(new_n701_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n738_), .A2(G36gat), .A3(new_n672_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(KEYINPUT46), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n737_), .B(new_n741_), .C1(new_n743_), .C2(KEYINPUT46), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1329gat));
  NAND4_X1  g546(.A1(new_n726_), .A2(new_n732_), .A3(G43gat), .A4(new_n613_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n478_), .B1(new_n738_), .B2(new_n612_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(G1330gat));
  OR3_X1    g551(.A1(new_n738_), .A2(G50gat), .A3(new_n408_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n726_), .A2(new_n732_), .A3(new_n407_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n754_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT109), .B1(new_n754_), .B2(G50gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(G1331gat));
  NAND3_X1  g556(.A1(new_n336_), .A2(new_n339_), .A3(new_n312_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n663_), .B(new_n759_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n761_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n762_), .A2(G57gat), .A3(new_n624_), .A4(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n765_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n663_), .A2(new_n714_), .A3(new_n335_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n314_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G57gat), .B1(new_n770_), .B2(new_n624_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n766_), .A2(new_n767_), .A3(new_n771_), .ZN(G1332gat));
  OR3_X1    g571(.A1(new_n769_), .A2(G64gat), .A3(new_n672_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n762_), .A2(new_n676_), .A3(new_n763_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G64gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G64gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(G1333gat));
  NAND3_X1  g577(.A1(new_n762_), .A2(new_n613_), .A3(new_n763_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(G71gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G71gat), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n613_), .A2(new_n472_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT112), .ZN(new_n784_));
  OAI22_X1  g583(.A1(new_n781_), .A2(new_n782_), .B1(new_n769_), .B2(new_n784_), .ZN(G1334gat));
  OR3_X1    g584(.A1(new_n769_), .A2(G78gat), .A3(new_n408_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n762_), .A2(new_n407_), .A3(new_n763_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(new_n788_), .A3(G78gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n787_), .B2(G78gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(G1335gat));
  NOR3_X1   g590(.A1(new_n260_), .A2(new_n337_), .A3(new_n312_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n708_), .A2(new_n717_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n721_), .A2(new_n722_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G85gat), .B1(new_n797_), .B2(new_n539_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n768_), .A2(new_n699_), .ZN(new_n799_));
  OR3_X1    g598(.A1(new_n799_), .A2(G85gat), .A3(new_n539_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1336gat));
  OAI21_X1  g600(.A(G92gat), .B1(new_n797_), .B2(new_n672_), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n799_), .A2(G92gat), .A3(new_n672_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1337gat));
  AND4_X1   g603(.A1(new_n613_), .A2(new_n768_), .A3(new_n211_), .A4(new_n699_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(KEYINPUT113), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n797_), .A2(new_n612_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n470_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI211_X1 g608(.A(KEYINPUT52), .B(new_n212_), .C1(new_n796_), .C2(new_n407_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n731_), .A2(new_n407_), .A3(new_n792_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(G106gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n407_), .A2(new_n212_), .ZN(new_n814_));
  OAI22_X1  g613(.A1(new_n810_), .A2(new_n813_), .B1(new_n799_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT53), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817_));
  OAI221_X1 g616(.A(new_n817_), .B1(new_n799_), .B2(new_n814_), .C1(new_n810_), .C2(new_n813_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1339gat));
  NOR2_X1   g618(.A1(new_n676_), .A2(new_n407_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n612_), .A2(new_n539_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n236_), .A2(new_n243_), .A3(new_n238_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n241_), .A2(KEYINPUT55), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n243_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n252_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n828_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n337_), .A2(new_n253_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n828_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(KEYINPUT116), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n251_), .A2(new_n253_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n323_), .A2(new_n324_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n328_), .A2(new_n329_), .A3(new_n325_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n321_), .A3(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT117), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n331_), .A2(new_n321_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n834_), .A2(new_n837_), .B1(new_n838_), .B2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT118), .B(new_n823_), .C1(new_n845_), .C2(new_n284_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n834_), .A2(new_n837_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n838_), .A2(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT57), .A3(new_n698_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n831_), .A2(new_n833_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n844_), .A2(new_n253_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n851_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n852_), .A2(KEYINPUT58), .A3(new_n253_), .A4(new_n844_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n290_), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n846_), .A2(new_n850_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n849_), .B2(new_n698_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(KEYINPUT118), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n313_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n759_), .A2(KEYINPUT114), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n255_), .A2(new_n256_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n758_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n862_), .A2(new_n863_), .A3(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OR3_X1    g667(.A1(new_n866_), .A2(new_n290_), .A3(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n866_), .B2(new_n290_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n822_), .B1(new_n861_), .B2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n420_), .A3(new_n337_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n822_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT59), .B1(new_n874_), .B2(KEYINPUT120), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(KEYINPUT120), .B2(new_n874_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n856_), .A2(new_n290_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n854_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(KEYINPUT58), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n877_), .B1(new_n859_), .B2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n845_), .A2(new_n284_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n857_), .B(KEYINPUT121), .C1(new_n883_), .C2(KEYINPUT57), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(new_n884_), .A3(new_n850_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n313_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n876_), .B1(new_n886_), .B2(new_n871_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n872_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n869_), .A2(new_n870_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n883_), .B2(KEYINPUT57), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n893_), .A2(new_n857_), .A3(new_n850_), .A4(new_n846_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n891_), .B1(new_n894_), .B2(new_n313_), .ZN(new_n895_));
  OAI211_X1 g694(.A(KEYINPUT119), .B(KEYINPUT59), .C1(new_n895_), .C2(new_n822_), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n340_), .B(new_n887_), .C1(new_n890_), .C2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n873_), .B1(new_n897_), .B2(new_n420_), .ZN(G1340gat));
  OAI21_X1  g697(.A(new_n418_), .B1(new_n260_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n872_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n418_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n260_), .B(new_n887_), .C1(new_n890_), .C2(new_n896_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n418_), .ZN(G1341gat));
  NAND3_X1  g701(.A1(new_n872_), .A2(new_n415_), .A3(new_n312_), .ZN(new_n903_));
  AOI211_X1 g702(.A(new_n313_), .B(new_n887_), .C1(new_n890_), .C2(new_n896_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n415_), .ZN(G1342gat));
  AOI211_X1 g704(.A(new_n698_), .B(new_n822_), .C1(new_n861_), .C2(new_n871_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT122), .B1(new_n906_), .B2(G134gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n872_), .A2(new_n284_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(new_n909_), .A3(new_n413_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n887_), .B1(new_n890_), .B2(new_n896_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n705_), .A2(new_n413_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1343gat));
  NOR3_X1   g713(.A1(new_n613_), .A2(new_n408_), .A3(new_n539_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n672_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n895_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n337_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n663_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(new_n922_), .A3(new_n312_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n861_), .A2(new_n871_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n924_), .A2(new_n672_), .A3(new_n312_), .A4(new_n915_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT123), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT61), .B(G155gat), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n923_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n923_), .B2(new_n926_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1346gat));
  INV_X1    g729(.A(new_n917_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G162gat), .B1(new_n931_), .B2(new_n705_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n917_), .A2(new_n355_), .A3(new_n284_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1347gat));
  NAND2_X1  g733(.A1(new_n886_), .A2(new_n871_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n672_), .A2(new_n612_), .A3(new_n624_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT124), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n407_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n935_), .A2(new_n337_), .A3(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(G169gat), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n940_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n944_));
  INV_X1    g743(.A(new_n542_), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n943_), .B(new_n944_), .C1(new_n945_), .C2(new_n940_), .ZN(G1348gat));
  NAND2_X1  g745(.A1(new_n935_), .A2(new_n939_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n663_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n895_), .A2(new_n407_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n938_), .A2(new_n444_), .A3(new_n260_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n949_), .A2(new_n458_), .B1(new_n950_), .B2(new_n951_), .ZN(G1349gat));
  NOR3_X1   g751(.A1(new_n947_), .A2(new_n557_), .A3(new_n313_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n950_), .A2(new_n312_), .A3(new_n937_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n434_), .B2(new_n954_), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n947_), .B2(new_n705_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n284_), .A2(new_n558_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n947_), .B2(new_n957_), .ZN(G1351gat));
  NOR3_X1   g757(.A1(new_n672_), .A2(new_n613_), .A3(new_n618_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  OAI21_X1  g759(.A(KEYINPUT125), .B1(new_n895_), .B2(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n924_), .A2(new_n962_), .A3(new_n959_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n963_), .ZN(new_n964_));
  AND3_X1   g763(.A1(new_n964_), .A2(G197gat), .A3(new_n337_), .ZN(new_n965_));
  AOI21_X1  g764(.A(G197gat), .B1(new_n964_), .B2(new_n337_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1352gat));
  AOI21_X1  g766(.A(new_n260_), .B1(new_n961_), .B2(new_n963_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(new_n970_));
  XOR2_X1   g769(.A(KEYINPUT126), .B(G204gat), .Z(new_n971_));
  OAI21_X1  g770(.A(new_n970_), .B1(new_n968_), .B2(new_n971_), .ZN(G1353gat));
  XNOR2_X1  g771(.A(KEYINPUT63), .B(G211gat), .ZN(new_n973_));
  AOI211_X1 g772(.A(new_n313_), .B(new_n973_), .C1(new_n961_), .C2(new_n963_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n964_), .A2(new_n312_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n974_), .B1(new_n975_), .B2(new_n976_), .ZN(G1354gat));
  INV_X1    g776(.A(G218gat), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n964_), .A2(new_n978_), .A3(new_n284_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n705_), .B1(new_n961_), .B2(new_n963_), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n979_), .B1(new_n980_), .B2(new_n978_), .ZN(G1355gat));
endmodule


