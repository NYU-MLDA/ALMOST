//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G183gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT83), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT83), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G183gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n203_), .B1(new_n209_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n212_), .A2(new_n213_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT84), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT84), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n216_), .B(new_n217_), .C1(new_n223_), .C2(KEYINPUT24), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT24), .B1(new_n221_), .B2(new_n222_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT86), .B1(new_n225_), .B2(new_n214_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n228_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(G169gat), .B2(G176gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT85), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n234_), .A2(new_n221_), .A3(new_n237_), .A4(new_n222_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n232_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n215_), .B1(new_n227_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G71gat), .B(G99gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G43gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n240_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(G15gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT30), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT31), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n247_), .A2(new_n254_), .A3(new_n248_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G204gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT92), .B1(new_n259_), .B2(G197gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261_));
  INV_X1    g060(.A(G197gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(G204gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT92), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(new_n262_), .A3(G204gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n259_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n260_), .A2(new_n263_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT21), .ZN(new_n268_));
  INV_X1    g067(.A(G218gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G211gat), .ZN(new_n270_));
  INV_X1    g069(.A(G211gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G218gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n268_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G211gat), .B(G218gat), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n275_), .A2(new_n278_), .A3(new_n274_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n240_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT19), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n279_), .B1(new_n268_), .B2(new_n276_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n229_), .A2(new_n204_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n287_), .A2(KEYINPUT96), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT96), .B1(new_n287_), .B2(new_n288_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n228_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n225_), .A2(new_n214_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(new_n235_), .ZN(new_n293_));
  OR2_X1    g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n217_), .A2(new_n294_), .B1(G169gat), .B2(G176gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n219_), .A2(KEYINPUT22), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT22), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G169gat), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n296_), .A2(new_n298_), .A3(KEYINPUT97), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT97), .B1(new_n296_), .B2(new_n298_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n220_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n295_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n286_), .A2(new_n293_), .A3(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n282_), .A2(KEYINPUT20), .A3(new_n285_), .A4(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n293_), .A2(new_n302_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n281_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n286_), .B(new_n215_), .C1(new_n227_), .C2(new_n239_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT20), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT98), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n284_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n309_), .B1(new_n308_), .B2(new_n284_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n304_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G8gat), .B(G36gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n317_), .B(new_n304_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT27), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(KEYINPUT87), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n324_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n322_), .A2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n323_), .A2(KEYINPUT1), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n340_), .B1(new_n341_), .B2(new_n322_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n325_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n343_), .A2(new_n328_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(new_n246_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G85gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT0), .B(G57gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n246_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n346_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n325_), .A2(new_n326_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n358_), .A2(new_n331_), .A3(new_n335_), .A4(new_n336_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n359_), .A2(new_n324_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n246_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n361_), .A3(KEYINPUT4), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n360_), .A2(KEYINPUT4), .A3(new_n246_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n350_), .B(new_n355_), .C1(new_n364_), .C2(new_n348_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n348_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n347_), .A2(new_n349_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n354_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G22gat), .B(G50gat), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n360_), .B2(new_n373_), .ZN(new_n374_));
  AND4_X1   g173(.A1(new_n373_), .A2(new_n338_), .A3(new_n345_), .A4(new_n372_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n371_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n372_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n346_), .B2(KEYINPUT29), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n360_), .A2(new_n373_), .A3(new_n372_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n370_), .A3(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(KEYINPUT94), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT95), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT95), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n376_), .A2(new_n380_), .A3(KEYINPUT94), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT94), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n374_), .A2(new_n375_), .A3(new_n371_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n370_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(G228gat), .B1(KEYINPUT90), .B2(G233gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(KEYINPUT90), .B2(G233gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n281_), .B2(KEYINPUT89), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT93), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n281_), .B(new_n394_), .C1(new_n373_), .C2(new_n360_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n373_), .B1(new_n338_), .B2(new_n345_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n396_), .B1(new_n397_), .B2(new_n286_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n392_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n392_), .A3(new_n398_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n389_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n385_), .A2(new_n402_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n395_), .A2(new_n392_), .A3(new_n398_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(new_n399_), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n389_), .A2(new_n405_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n369_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n305_), .A2(KEYINPUT101), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT101), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n293_), .A2(new_n302_), .A3(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n286_), .A3(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n240_), .B2(new_n281_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n285_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n308_), .A2(new_n284_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n318_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n320_), .A2(KEYINPUT27), .A3(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n321_), .A2(new_n407_), .A3(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n385_), .B(new_n402_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n357_), .A2(new_n361_), .A3(new_n349_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n355_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n364_), .B2(new_n348_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n368_), .A2(KEYINPUT33), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n424_), .B(new_n354_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(new_n320_), .A3(new_n319_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n317_), .A2(KEYINPUT32), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT102), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n365_), .A2(new_n368_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n304_), .B(new_n428_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n434_));
  OAI211_X1 g233(.A(KEYINPUT102), .B(new_n429_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n419_), .B1(new_n427_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n258_), .B1(new_n418_), .B2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n321_), .A2(new_n417_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n419_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n258_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n439_), .A2(new_n369_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G29gat), .B(G36gat), .Z(new_n444_));
  XOR2_X1   g243(.A(G43gat), .B(G50gat), .Z(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G1gat), .ZN(new_n447_));
  INV_X1    g246(.A(G8gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT14), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT78), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(KEYINPUT78), .B(KEYINPUT14), .C1(new_n447_), .C2(new_n448_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G15gat), .B(G22gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT79), .ZN(new_n455_));
  XOR2_X1   g254(.A(G1gat), .B(G8gat), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n455_), .A2(new_n457_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n446_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n455_), .A2(new_n457_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n446_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n458_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G229gat), .A3(G233gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT80), .Z(new_n468_));
  NAND2_X1  g267(.A1(new_n462_), .A2(new_n458_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n446_), .B(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n461_), .B(new_n468_), .C1(new_n469_), .C2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G113gat), .B(G141gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT81), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT82), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G169gat), .B(G197gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n466_), .A2(new_n472_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n466_), .B2(new_n472_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n443_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT103), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n443_), .A2(KEYINPUT103), .A3(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT77), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(KEYINPUT66), .ZN(new_n492_));
  INV_X1    g291(.A(G99gat), .ZN(new_n493_));
  INV_X1    g292(.A(G106gat), .ZN(new_n494_));
  OAI22_X1  g293(.A1(new_n490_), .A2(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(KEYINPUT66), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n497_));
  AND2_X1   g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT10), .B(G99gat), .ZN(new_n501_));
  AND2_X1   g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT9), .ZN(new_n503_));
  NOR2_X1   g302(.A1(G85gat), .A2(G92gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n503_), .B1(new_n504_), .B2(KEYINPUT65), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(KEYINPUT65), .B2(new_n503_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT64), .B(G92gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT9), .B1(new_n507_), .B2(G85gat), .ZN(new_n508_));
  OAI221_X1 g307(.A(new_n500_), .B1(G106gat), .B2(new_n501_), .C1(new_n506_), .C2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n502_), .A2(new_n504_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT8), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n498_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(G99gat), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n494_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n493_), .A2(new_n494_), .A3(KEYINPUT67), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT7), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT68), .B1(new_n515_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT68), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n500_), .A2(new_n524_), .A3(new_n521_), .A4(new_n519_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n512_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n518_), .B1(new_n517_), .B2(new_n494_), .ZN(new_n527_));
  NOR4_X1   g326(.A1(new_n516_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT69), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT69), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n519_), .A2(new_n521_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n500_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n511_), .B1(new_n532_), .B2(new_n510_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n509_), .B1(new_n526_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n446_), .B(KEYINPUT15), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n446_), .B(new_n509_), .C1(new_n526_), .C2(new_n533_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT34), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT74), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n536_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G190gat), .B(G218gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT73), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n542_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n544_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n537_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n545_), .A2(KEYINPUT75), .A3(new_n551_), .A4(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n556_), .A2(KEYINPUT37), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n549_), .B(KEYINPUT36), .ZN(new_n558_));
  AND4_X1   g357(.A1(new_n554_), .A2(new_n536_), .A3(new_n537_), .A4(new_n542_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n554_), .B1(new_n553_), .B2(new_n537_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n545_), .A2(new_n551_), .A3(new_n555_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT75), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(new_n562_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT76), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT76), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n561_), .A2(new_n562_), .A3(new_n568_), .A4(new_n565_), .ZN(new_n569_));
  AOI221_X4 g368(.A(new_n488_), .B1(new_n557_), .B2(new_n564_), .C1(new_n567_), .C2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n569_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n557_), .A2(new_n564_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT77), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G57gat), .B(G64gat), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT11), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT11), .ZN(new_n577_));
  XOR2_X1   g376(.A(G71gat), .B(G78gat), .Z(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n534_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n509_), .B(new_n581_), .C1(new_n526_), .C2(new_n533_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(KEYINPUT12), .A3(new_n584_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n534_), .A2(new_n590_), .A3(new_n582_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n586_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G120gat), .B(G148gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT5), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n593_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n586_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n587_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT70), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n599_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(KEYINPUT70), .B(new_n597_), .C1(new_n587_), .C2(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT71), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT13), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n606_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n604_), .A2(new_n607_), .A3(new_n608_), .A4(new_n605_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n581_), .B(new_n614_), .Z(new_n615_));
  XNOR2_X1  g414(.A(new_n469_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT17), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT16), .ZN(new_n619_));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n616_), .A2(new_n617_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(KEYINPUT17), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n616_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n574_), .A2(new_n613_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n487_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT104), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n433_), .A2(new_n447_), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n561_), .A2(new_n562_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n626_), .B(new_n634_), .C1(new_n438_), .C2(new_n442_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n613_), .A2(new_n481_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n637_), .B2(new_n369_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n630_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n632_), .A2(new_n638_), .A3(new_n639_), .ZN(G1324gat));
  OAI21_X1  g439(.A(G8gat), .B1(new_n637_), .B2(new_n439_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT39), .ZN(new_n642_));
  INV_X1    g441(.A(new_n439_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n448_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n629_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n642_), .B(new_n646_), .C1(new_n629_), .C2(new_n644_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n637_), .B2(new_n258_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n652_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n628_), .A2(G15gat), .A3(new_n258_), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(G1326gat));
  OAI21_X1  g458(.A(G22gat), .B1(new_n637_), .B2(new_n440_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n440_), .A2(G22gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n628_), .B2(new_n662_), .ZN(G1327gat));
  AND2_X1   g462(.A1(new_n611_), .A2(new_n612_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n625_), .A2(new_n633_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G29gat), .B1(new_n667_), .B2(new_n433_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n571_), .A2(new_n572_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n488_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n571_), .A2(KEYINPUT77), .A3(new_n572_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n443_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n673_), .A3(new_n671_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(KEYINPUT43), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n574_), .B(new_n443_), .C1(new_n673_), .C2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n664_), .A2(new_n482_), .A3(new_n626_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT44), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n682_), .B(new_n679_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n433_), .A2(G29gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n668_), .B1(new_n684_), .B2(new_n685_), .ZN(G1328gat));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  INV_X1    g486(.A(G36gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n684_), .B2(new_n643_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n439_), .A2(G36gat), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n667_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n667_), .B2(new_n691_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n687_), .B1(new_n689_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n694_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n681_), .A2(new_n683_), .A3(new_n439_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n696_), .B(KEYINPUT46), .C1(new_n697_), .C2(new_n688_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(G1329gat));
  NAND3_X1  g498(.A1(new_n684_), .A2(G43gat), .A3(new_n441_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n667_), .A2(new_n441_), .ZN(new_n703_));
  INV_X1    g502(.A(G43gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  AOI211_X1 g504(.A(KEYINPUT109), .B(G43gat), .C1(new_n667_), .C2(new_n441_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n700_), .B(new_n701_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n441_), .A2(G43gat), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n681_), .A2(new_n683_), .A3(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT47), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n667_), .B2(new_n419_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n419_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n684_), .B2(new_n714_), .ZN(G1331gat));
  NOR2_X1   g514(.A1(new_n574_), .A2(new_n626_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n482_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(new_n443_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G57gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n433_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n635_), .A2(new_n717_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n369_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1332gat));
  NOR2_X1   g522(.A1(new_n439_), .A2(G64gat), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT112), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n718_), .A2(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G64gat), .B1(new_n721_), .B2(new_n439_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT111), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(G64gat), .C1(new_n721_), .C2(new_n439_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n728_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n728_), .B2(new_n730_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n726_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT113), .B(new_n726_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n721_), .B2(new_n258_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n258_), .A2(G71gat), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT115), .Z(new_n743_));
  NAND2_X1  g542(.A1(new_n718_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n721_), .B2(new_n440_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT50), .ZN(new_n747_));
  INV_X1    g546(.A(G78gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n718_), .A2(new_n748_), .A3(new_n419_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1335gat));
  AND3_X1   g549(.A1(new_n717_), .A2(new_n443_), .A3(new_n665_), .ZN(new_n751_));
  INV_X1    g550(.A(G85gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n433_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n717_), .A2(new_n626_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT117), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n717_), .A2(KEYINPUT117), .A3(new_n626_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n678_), .B2(KEYINPUT116), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n759_), .A2(new_n369_), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n753_), .B1(new_n762_), .B2(new_n752_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT118), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT118), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n753_), .C1(new_n762_), .C2(new_n752_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1336gat));
  AOI21_X1  g566(.A(G92gat), .B1(new_n751_), .B2(new_n643_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n759_), .A2(new_n761_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n643_), .A2(new_n507_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(G1337gat));
  INV_X1    g570(.A(new_n501_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n751_), .A2(new_n441_), .A3(new_n772_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n759_), .A2(new_n258_), .A3(new_n761_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n493_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT51), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n773_), .C1(new_n774_), .C2(new_n493_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n678_), .A2(new_n758_), .A3(new_n419_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G106gat), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n751_), .A2(new_n494_), .A3(new_n419_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT119), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n784_), .A3(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n783_), .A2(new_n784_), .A3(new_n786_), .A4(new_n788_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n716_), .A2(new_n793_), .A3(new_n481_), .A4(new_n664_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n670_), .A2(new_n671_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n795_), .A2(new_n664_), .A3(new_n481_), .A4(new_n625_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT54), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n477_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n459_), .A2(new_n471_), .A3(new_n460_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n463_), .B1(new_n462_), .B2(new_n458_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT121), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n468_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n800_), .A2(new_n801_), .A3(KEYINPUT121), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n799_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n806_), .A2(new_n478_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n604_), .A2(new_n807_), .A3(new_n605_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT122), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n589_), .A2(new_n600_), .A3(new_n591_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n593_), .A2(KEYINPUT55), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n598_), .B1(new_n601_), .B2(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n814_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n482_), .B(new_n599_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n604_), .A2(new_n807_), .A3(KEYINPUT122), .A4(new_n605_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n810_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(KEYINPUT57), .A3(new_n633_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n599_), .A2(new_n478_), .A3(new_n806_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n821_), .B(KEYINPUT58), .C1(new_n815_), .C2(new_n816_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n670_), .A2(new_n824_), .A3(new_n671_), .A4(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n819_), .B2(new_n633_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n626_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n798_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n643_), .A2(new_n419_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n433_), .A3(new_n441_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n831_), .A2(new_n832_), .A3(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n820_), .B(new_n826_), .C1(new_n829_), .C2(KEYINPUT124), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n829_), .A2(KEYINPUT124), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n626_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n834_), .B1(new_n839_), .B2(new_n798_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n836_), .B(new_n482_), .C1(new_n840_), .C2(new_n832_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G113gat), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n843_), .A3(new_n482_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1340gat));
  OAI211_X1 g644(.A(new_n836_), .B(new_n613_), .C1(new_n840_), .C2(new_n832_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G120gat), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n664_), .A2(KEYINPUT60), .ZN(new_n848_));
  MUX2_X1   g647(.A(new_n848_), .B(KEYINPUT60), .S(G120gat), .Z(new_n849_));
  NAND2_X1  g648(.A1(new_n840_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(G1341gat));
  NAND2_X1  g650(.A1(new_n625_), .A2(G127gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT125), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n836_), .B(new_n853_), .C1(new_n840_), .C2(new_n832_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G127gat), .B1(new_n840_), .B2(new_n625_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1342gat));
  OAI211_X1 g656(.A(new_n836_), .B(new_n574_), .C1(new_n840_), .C2(new_n832_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G134gat), .ZN(new_n859_));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n840_), .A2(new_n860_), .A3(new_n634_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1343gat));
  NAND2_X1  g661(.A1(new_n839_), .A2(new_n798_), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n643_), .A2(new_n369_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n482_), .A3(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n613_), .A3(new_n864_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g667(.A1(new_n863_), .A2(new_n625_), .A3(new_n864_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  INV_X1    g670(.A(G162gat), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n863_), .A2(new_n872_), .A3(new_n634_), .A4(new_n864_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n863_), .A2(new_n574_), .A3(new_n864_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n872_), .ZN(G1347gat));
  NOR3_X1   g674(.A1(new_n439_), .A2(new_n433_), .A3(new_n258_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n440_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n798_), .B2(new_n830_), .ZN(new_n878_));
  AOI211_X1 g677(.A(KEYINPUT62), .B(new_n219_), .C1(new_n878_), .C2(new_n482_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n482_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(G169gat), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n878_), .B(new_n482_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n882_), .B2(new_n883_), .ZN(G1348gat));
  AOI211_X1 g683(.A(new_n664_), .B(new_n877_), .C1(new_n798_), .C2(new_n830_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT126), .B1(new_n885_), .B2(G176gat), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n887_));
  INV_X1    g686(.A(new_n877_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n831_), .A2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n887_), .B(new_n220_), .C1(new_n889_), .C2(new_n664_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n419_), .B1(new_n839_), .B2(new_n798_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n613_), .A2(G176gat), .A3(new_n876_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n886_), .A2(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n625_), .A3(new_n876_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n208_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n626_), .A2(new_n290_), .A3(new_n289_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n894_), .A2(new_n895_), .B1(new_n878_), .B2(new_n896_), .ZN(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n889_), .B2(new_n795_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n878_), .A2(new_n228_), .A3(new_n634_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1351gat));
  NOR3_X1   g699(.A1(new_n439_), .A2(new_n407_), .A3(new_n441_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n839_), .B2(new_n798_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n482_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n613_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n908_), .A2(new_n271_), .A3(KEYINPUT127), .ZN(new_n909_));
  AOI211_X1 g708(.A(new_n909_), .B(new_n626_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n903_), .A2(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(KEYINPUT127), .B1(new_n908_), .B2(new_n271_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1354gat));
  INV_X1    g712(.A(new_n903_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G218gat), .B1(new_n914_), .B2(new_n795_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n903_), .A2(new_n269_), .A3(new_n634_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1355gat));
endmodule


