//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT74), .B(G15gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(G22gat), .ZN(new_n209_));
  INV_X1    g008(.A(G1gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n214_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n207_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n219_));
  INV_X1    g018(.A(new_n206_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n206_), .A2(new_n215_), .A3(KEYINPUT76), .A4(new_n216_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n218_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n217_), .A2(new_n220_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n227_), .B2(new_n224_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G141gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT77), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G169gat), .B(G197gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n230_), .B(new_n231_), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n232_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n225_), .B(new_n234_), .C1(new_n227_), .C2(new_n224_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n235_), .A2(KEYINPUT78), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(KEYINPUT78), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n233_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G141gat), .B(G148gat), .Z(new_n239_));
  NAND2_X1  g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT1), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT83), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n245_), .A2(KEYINPUT84), .A3(G155gat), .A4(G162gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT82), .ZN(new_n248_));
  INV_X1    g047(.A(G155gat), .ZN(new_n249_));
  INV_X1    g048(.A(G162gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n240_), .A2(KEYINPUT1), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n251_), .B(new_n252_), .C1(new_n253_), .C2(KEYINPUT84), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n239_), .B1(new_n247_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT85), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT2), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT2), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(KEYINPUT85), .A3(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n261_));
  OR3_X1    g060(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n258_), .A2(new_n260_), .A3(new_n261_), .A4(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n251_), .A2(new_n240_), .A3(new_n252_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n255_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G113gat), .B(G120gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n270_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G225gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(KEYINPUT4), .A3(new_n272_), .ZN(new_n277_));
  OR3_X1    g076(.A1(new_n267_), .A2(KEYINPUT4), .A3(new_n270_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n274_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G85gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G57gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  OR3_X1    g082(.A1(new_n276_), .A2(new_n279_), .A3(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n283_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G228gat), .ZN(new_n288_));
  INV_X1    g087(.A(G233gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT91), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT91), .B1(new_n288_), .B2(new_n289_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G197gat), .B(G204gat), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT90), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(KEYINPUT90), .ZN(new_n296_));
  INV_X1    g095(.A(G218gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G211gat), .ZN(new_n298_));
  INV_X1    g097(.A(G211gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G218gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n295_), .A2(new_n296_), .A3(KEYINPUT21), .A4(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(G197gat), .A2(G204gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G197gat), .A2(G204gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n301_), .B1(KEYINPUT21), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT21), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT88), .B1(new_n294_), .B2(new_n308_), .ZN(new_n309_));
  OAI211_X1 g108(.A(KEYINPUT88), .B(new_n308_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n307_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT89), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n306_), .B2(KEYINPUT21), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n310_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(KEYINPUT89), .A3(new_n307_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n303_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n255_), .B2(new_n265_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n292_), .B(new_n293_), .C1(new_n319_), .C2(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n317_), .A2(KEYINPUT89), .A3(new_n307_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT89), .B1(new_n317_), .B2(new_n307_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n302_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n321_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n325_), .A2(new_n291_), .A3(new_n290_), .A4(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n322_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n328_), .B1(new_n322_), .B2(new_n327_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n255_), .A2(new_n320_), .A3(new_n265_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT86), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT28), .B(G22gat), .ZN(new_n333_));
  INV_X1    g132(.A(G50gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT86), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n255_), .A2(new_n265_), .A3(new_n336_), .A4(new_n320_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n332_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n339_), .A2(new_n340_), .A3(KEYINPUT87), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n332_), .A2(new_n337_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n335_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n342_), .B1(new_n345_), .B2(new_n338_), .ZN(new_n346_));
  OAI22_X1  g145(.A1(new_n329_), .A2(new_n330_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n322_), .A2(new_n327_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n328_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n322_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n345_), .A2(new_n338_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n347_), .A2(KEYINPUT92), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT93), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT92), .ZN(new_n356_));
  OAI221_X1 g155(.A(new_n356_), .B1(new_n341_), .B2(new_n346_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n355_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n287_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT27), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT25), .B(G183gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT23), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(G183gat), .A3(G190gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n364_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT79), .ZN(new_n375_));
  INV_X1    g174(.A(new_n370_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(KEYINPUT24), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G169gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT22), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G169gat), .ZN(new_n381_));
  INV_X1    g180(.A(G176gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n375_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n368_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G183gat), .ZN(new_n387_));
  INV_X1    g186(.A(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n366_), .A2(new_n368_), .A3(new_n385_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n373_), .A2(new_n377_), .B1(new_n384_), .B2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n392_), .B(new_n302_), .C1(new_n323_), .C2(new_n324_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n376_), .A2(new_n374_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n370_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n396_), .A2(new_n364_), .A3(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n386_), .A2(new_n390_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n369_), .A2(new_n389_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n398_), .A2(new_n399_), .B1(new_n384_), .B2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n393_), .B(KEYINPUT20), .C1(new_n319_), .C2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT19), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT18), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n407_), .B(new_n408_), .Z(new_n409_));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n319_), .B2(new_n401_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n404_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n392_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n325_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n405_), .A2(new_n409_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n409_), .B1(new_n405_), .B2(new_n415_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n361_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT96), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT96), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(new_n361_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n405_), .A2(new_n409_), .A3(new_n415_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT95), .ZN(new_n424_));
  INV_X1    g223(.A(new_n409_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n402_), .A2(new_n404_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n412_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n424_), .A2(KEYINPUT27), .A3(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n423_), .A2(KEYINPUT95), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n422_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT97), .B1(new_n360_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n354_), .A2(new_n357_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT93), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n419_), .A2(new_n421_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .A4(new_n287_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n285_), .B(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n283_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n277_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OR3_X1    g244(.A1(new_n445_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n409_), .A2(KEYINPUT32), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n405_), .A2(new_n415_), .A3(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n426_), .A2(new_n427_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(new_n447_), .ZN(new_n450_));
  OAI22_X1  g249(.A1(new_n442_), .A2(new_n446_), .B1(new_n287_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n433_), .A2(new_n440_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT98), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G71gat), .B(G99gat), .ZN(new_n455_));
  INV_X1    g254(.A(G43gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n392_), .B(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G227gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G15gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT30), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(new_n270_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n464_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n453_), .A2(new_n454_), .A3(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n437_), .A2(new_n432_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n468_), .A2(new_n286_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n454_), .B1(new_n453_), .B2(new_n468_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n238_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT99), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n453_), .A2(new_n468_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT98), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n472_), .A3(new_n469_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT99), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n238_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G232gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT34), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT35), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AOI211_X1 g286(.A(G99gat), .B(G106gat), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(KEYINPUT65), .B2(KEYINPUT7), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT6), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n489_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G85gat), .B(G92gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT8), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT9), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(G85gat), .A3(G92gat), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n494_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT10), .B(G99gat), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI221_X1 g304(.A(new_n503_), .B1(new_n501_), .B2(new_n496_), .C1(G106gat), .C2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n500_), .A2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n207_), .A2(KEYINPUT71), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT71), .B1(new_n207_), .B2(new_n507_), .ZN(new_n509_));
  OAI221_X1 g308(.A(new_n487_), .B1(new_n220_), .B2(new_n507_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n485_), .A2(new_n486_), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  XOR2_X1   g311(.A(G190gat), .B(G218gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(G134gat), .B(G162gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT72), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n510_), .A2(new_n511_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n510_), .A2(new_n511_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n515_), .B(KEYINPUT36), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n519_), .A2(new_n524_), .A3(KEYINPUT37), .ZN(new_n525_));
  INV_X1    g324(.A(new_n523_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n522_), .B2(KEYINPUT73), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n520_), .A2(new_n528_), .A3(new_n521_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n527_), .A2(new_n529_), .B1(new_n512_), .B2(new_n518_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n525_), .B1(new_n530_), .B2(KEYINPUT37), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n217_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT11), .Z(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT67), .B(G71gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(G78gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n538_), .B1(new_n539_), .B2(new_n537_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n533_), .B(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G127gat), .B(G155gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT16), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G183gat), .B(G211gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n542_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT75), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n546_), .A2(new_n547_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n542_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n540_), .B1(new_n500_), .B2(new_n506_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n500_), .A2(new_n506_), .A3(new_n540_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(KEYINPUT68), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(G230gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(new_n289_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n558_), .B(new_n560_), .C1(KEYINPUT68), .C2(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(KEYINPUT12), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(new_n555_), .ZN(new_n563_));
  AOI211_X1 g362(.A(KEYINPUT12), .B(new_n540_), .C1(new_n500_), .C2(new_n506_), .ZN(new_n564_));
  OAI22_X1  g363(.A1(new_n563_), .A2(new_n564_), .B1(new_n559_), .B2(new_n289_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT5), .ZN(new_n568_));
  XOR2_X1   g367(.A(G176gat), .B(G204gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n570_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n571_), .A2(KEYINPUT13), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT13), .B1(new_n571_), .B2(new_n572_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n531_), .A2(new_n554_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n482_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT100), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n482_), .A2(KEYINPUT100), .A3(new_n577_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n287_), .A2(G1gat), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n580_), .A2(KEYINPUT38), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT101), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n238_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n576_), .A2(new_n586_), .A3(new_n554_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT102), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n527_), .A2(new_n529_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n519_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n479_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n588_), .B1(new_n479_), .B2(new_n590_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n587_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT103), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT103), .ZN(new_n596_));
  INV_X1    g395(.A(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n591_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n596_), .B1(new_n598_), .B2(new_n587_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n286_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n580_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n600_), .A2(G1gat), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n585_), .A2(new_n603_), .ZN(G1324gat));
  NAND4_X1  g403(.A1(new_n580_), .A2(new_n211_), .A3(new_n432_), .A4(new_n581_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n432_), .A3(new_n587_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n606_), .A2(new_n607_), .A3(G8gat), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n606_), .B2(G8gat), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT40), .B(new_n605_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(G1325gat));
  NAND2_X1  g413(.A1(new_n594_), .A2(KEYINPUT103), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n598_), .A2(new_n596_), .A3(new_n587_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n468_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT41), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(G15gat), .ZN(new_n620_));
  INV_X1    g419(.A(G15gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT41), .B1(new_n617_), .B2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n482_), .A2(new_n621_), .A3(new_n467_), .A4(new_n577_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT104), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n624_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n620_), .A2(new_n622_), .A3(new_n625_), .A4(new_n626_), .ZN(G1326gat));
  INV_X1    g426(.A(new_n437_), .ZN(new_n628_));
  OR3_X1    g427(.A1(new_n578_), .A2(G22gat), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n437_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(new_n631_), .A3(G22gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n630_), .B2(G22gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(G1327gat));
  NAND3_X1  g433(.A1(new_n530_), .A2(new_n554_), .A3(new_n575_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n476_), .B2(new_n481_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n286_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n575_), .A2(new_n238_), .A3(new_n554_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT43), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n531_), .B(new_n641_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n479_), .B2(new_n531_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT44), .B(new_n639_), .C1(new_n643_), .C2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT106), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n531_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n644_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n638_), .B1(new_n650_), .B2(new_n642_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n647_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n639_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n286_), .A2(G29gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n637_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  INV_X1    g459(.A(KEYINPUT108), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(KEYINPUT46), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n438_), .A2(G36gat), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n636_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n664_), .B1(new_n636_), .B2(new_n665_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n635_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n482_), .A2(new_n669_), .A3(new_n665_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT107), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n636_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(KEYINPUT45), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n668_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n438_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n654_), .B2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n662_), .B1(new_n674_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n650_), .A2(new_n642_), .ZN(new_n679_));
  AND4_X1   g478(.A1(new_n652_), .A2(new_n679_), .A3(KEYINPUT44), .A4(new_n639_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n652_), .B1(new_n651_), .B2(KEYINPUT44), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n676_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  INV_X1    g482(.A(new_n662_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n673_), .A4(new_n668_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n678_), .A2(new_n685_), .ZN(G1329gat));
  NOR2_X1   g485(.A1(new_n468_), .A2(new_n456_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n654_), .A2(new_n657_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n636_), .A2(new_n467_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n456_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT47), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(new_n693_), .A3(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1330gat));
  AOI21_X1  g494(.A(G50gat), .B1(new_n636_), .B2(new_n437_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n628_), .A2(new_n334_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n658_), .B2(new_n697_), .ZN(G1331gat));
  NAND3_X1  g497(.A1(new_n576_), .A2(new_n586_), .A3(new_n553_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n598_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G57gat), .B1(new_n287_), .B2(KEYINPUT109), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(KEYINPUT109), .B2(G57gat), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n479_), .A2(new_n586_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n531_), .A2(new_n554_), .A3(new_n575_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(new_n287_), .ZN(new_n707_));
  OAI22_X1  g506(.A1(new_n701_), .A2(new_n703_), .B1(new_n707_), .B2(G57gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT110), .ZN(G1332gat));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710_));
  INV_X1    g509(.A(new_n701_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n432_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n710_), .B1(new_n712_), .B2(G64gat), .ZN(new_n713_));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  AOI211_X1 g513(.A(KEYINPUT48), .B(new_n714_), .C1(new_n711_), .C2(new_n432_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n432_), .A2(new_n714_), .ZN(new_n716_));
  OAI22_X1  g515(.A1(new_n713_), .A2(new_n715_), .B1(new_n706_), .B2(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(KEYINPUT49), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n711_), .A2(new_n467_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G71gat), .ZN(new_n720_));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT49), .B(new_n721_), .C1(new_n711_), .C2(new_n467_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n467_), .A2(new_n721_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT111), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n720_), .A2(new_n722_), .B1(new_n706_), .B2(new_n724_), .ZN(G1334gat));
  OR3_X1    g524(.A1(new_n706_), .A2(G78gat), .A3(new_n628_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n437_), .B(new_n700_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G78gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G78gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT112), .ZN(G1335gat));
  NAND3_X1  g531(.A1(new_n576_), .A2(new_n586_), .A3(new_n554_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n679_), .A2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n287_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n590_), .A2(new_n553_), .A3(new_n575_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n704_), .A2(new_n737_), .ZN(new_n738_));
  OR3_X1    g537(.A1(new_n738_), .A2(G85gat), .A3(new_n287_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n735_), .B2(new_n438_), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n738_), .A2(G92gat), .A3(new_n438_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  NOR3_X1   g542(.A1(new_n738_), .A2(new_n468_), .A3(new_n505_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747_));
  INV_X1    g546(.A(G99gat), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n735_), .A2(new_n468_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n746_), .B(new_n747_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n744_), .B(KEYINPUT113), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n748_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT51), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n750_), .A2(new_n753_), .ZN(G1338gat));
  OR3_X1    g553(.A1(new_n738_), .A2(G106gat), .A3(new_n628_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n679_), .A2(new_n437_), .A3(new_n734_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n756_), .A2(G106gat), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n756_), .B2(G106gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n761_), .B(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n765_), .A2(KEYINPUT116), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n577_), .A2(new_n586_), .A3(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n519_), .A2(new_n524_), .A3(KEYINPUT37), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT37), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n590_), .B2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n771_), .A2(new_n586_), .A3(new_n553_), .A4(new_n575_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n768_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n556_), .A2(KEYINPUT12), .A3(new_n557_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n564_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n560_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT55), .B1(new_n778_), .B2(KEYINPUT117), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n565_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n777_), .A3(new_n560_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n779_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT56), .A3(new_n570_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT119), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n784_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n570_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n784_), .A2(new_n570_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n787_), .A2(new_n788_), .A3(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n236_), .A2(new_n237_), .ZN(new_n793_));
  AND4_X1   g592(.A1(G229gat), .A2(new_n218_), .A3(new_n223_), .A4(G233gat), .ZN(new_n794_));
  INV_X1    g593(.A(new_n227_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n234_), .B(new_n794_), .C1(new_n795_), .C2(new_n224_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n793_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(new_n571_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n792_), .A2(new_n798_), .A3(KEYINPUT58), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n531_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT120), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n801_), .A2(new_n531_), .A3(KEYINPUT120), .A4(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n238_), .A2(new_n571_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n791_), .B2(new_n785_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n571_), .A2(new_n572_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n797_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n811_), .A2(new_n530_), .B1(KEYINPUT118), .B2(KEYINPUT57), .ZN(new_n812_));
  NOR2_X1   g611(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n590_), .B(new_n813_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n805_), .A2(new_n806_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n775_), .B1(new_n554_), .B2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n470_), .A2(new_n467_), .A3(new_n286_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n768_), .A2(new_n774_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n553_), .B1(new_n815_), .B2(new_n803_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(KEYINPUT122), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n824_), .B(new_n553_), .C1(new_n815_), .C2(new_n803_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n818_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n828_));
  AND2_X1   g627(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI22_X1  g629(.A1(new_n819_), .A2(new_n820_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n586_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n819_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n586_), .A2(G113gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(G1340gat));
  OAI21_X1  g634(.A(G120gat), .B1(new_n831_), .B2(new_n575_), .ZN(new_n836_));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n575_), .B2(KEYINPUT60), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(KEYINPUT60), .B2(new_n837_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n836_), .B1(new_n833_), .B2(new_n839_), .ZN(G1341gat));
  OAI21_X1  g639(.A(G127gat), .B1(new_n831_), .B2(new_n554_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n554_), .A2(G127gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n833_), .B2(new_n842_), .ZN(G1342gat));
  OAI21_X1  g642(.A(G134gat), .B1(new_n831_), .B2(new_n771_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n590_), .A2(G134gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n833_), .B2(new_n845_), .ZN(G1343gat));
  NOR4_X1   g645(.A1(new_n628_), .A2(new_n432_), .A3(new_n467_), .A4(new_n287_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n817_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n238_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT123), .B(G141gat), .Z(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n576_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n816_), .A2(new_n554_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n553_), .B(new_n847_), .C1(new_n857_), .C2(new_n775_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT124), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(KEYINPUT124), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n856_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n861_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n859_), .A3(new_n855_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1346gat));
  OAI211_X1 g664(.A(new_n530_), .B(new_n847_), .C1(new_n857_), .C2(new_n775_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n250_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(KEYINPUT125), .A3(new_n250_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n771_), .A2(new_n250_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n869_), .A2(new_n870_), .B1(new_n849_), .B2(new_n871_), .ZN(G1347gat));
  NAND2_X1  g671(.A1(new_n432_), .A2(new_n471_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n437_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n238_), .B(new_n874_), .C1(new_n823_), .C2(new_n825_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n815_), .A2(new_n803_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n824_), .B1(new_n877_), .B2(new_n553_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n822_), .A2(KEYINPUT122), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n821_), .A3(new_n879_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n379_), .A2(new_n381_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n880_), .A2(new_n238_), .A3(new_n881_), .A4(new_n874_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT62), .B1(new_n875_), .B2(G169gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT126), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n875_), .A2(G169gat), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n882_), .A4(new_n876_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n885_), .A2(new_n890_), .ZN(G1348gat));
  NOR3_X1   g690(.A1(new_n826_), .A2(new_n437_), .A3(new_n873_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G176gat), .B1(new_n892_), .B2(new_n576_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n817_), .A2(new_n437_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n575_), .A2(new_n382_), .A3(new_n873_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  NAND4_X1  g695(.A1(new_n894_), .A2(new_n432_), .A3(new_n471_), .A4(new_n553_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n554_), .A2(new_n362_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n897_), .A2(new_n387_), .B1(new_n892_), .B2(new_n898_), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n363_), .A3(new_n530_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n892_), .A2(new_n531_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n902_), .B2(new_n388_), .ZN(G1351gat));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n360_), .A2(new_n467_), .A3(new_n438_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n817_), .B2(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n905_), .B(KEYINPUT127), .C1(new_n857_), .C2(new_n775_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n586_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(G197gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1352gat));
  AOI21_X1  g710(.A(new_n575_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n912_));
  INV_X1    g711(.A(G204gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1353gat));
  XNOR2_X1  g713(.A(KEYINPUT63), .B(G211gat), .ZN(new_n915_));
  AOI211_X1 g714(.A(new_n554_), .B(new_n915_), .C1(new_n907_), .C2(new_n908_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n907_), .A2(new_n908_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n553_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n916_), .B1(new_n918_), .B2(new_n919_), .ZN(G1354gat));
  NAND3_X1  g719(.A1(new_n917_), .A2(new_n297_), .A3(new_n530_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n771_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n297_), .B2(new_n922_), .ZN(G1355gat));
endmodule


