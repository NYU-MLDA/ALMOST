//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G71gat), .B(G78gat), .ZN(new_n205_));
  OR3_X1    g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n202_), .A2(new_n205_), .A3(KEYINPUT11), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(KEYINPUT79), .B(KEYINPUT14), .C1(new_n209_), .C2(new_n210_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G1gat), .B(G8gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n217_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n208_), .B(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G231gat), .A2(G233gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G127gat), .B(G155gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(G211gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT16), .B(G183gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n223_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(KEYINPUT17), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n223_), .A2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n232_), .B(KEYINPUT80), .Z(new_n233_));
  XNOR2_X1  g032(.A(G190gat), .B(G218gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G134gat), .B(G162gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT36), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(KEYINPUT76), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n237_), .A2(KEYINPUT76), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G232gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT34), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT35), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT6), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT6), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(G99gat), .A3(G106gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G85gat), .B(G92gat), .Z(new_n250_));
  AOI21_X1  g049(.A(new_n249_), .B1(KEYINPUT9), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT9), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(G85gat), .A3(G92gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT10), .B(G99gat), .Z(new_n254_));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n255_));
  INV_X1    g054(.A(G106gat), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n251_), .B(new_n253_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT65), .ZN(new_n260_));
  INV_X1    g059(.A(new_n250_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT7), .ZN(new_n262_));
  INV_X1    g061(.A(G99gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n256_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n264_), .A2(KEYINPUT68), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT68), .B1(new_n264_), .B2(new_n265_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n247_), .B1(G99gat), .B2(G106gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n245_), .A2(KEYINPUT6), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT67), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n261_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT8), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT69), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n278_));
  INV_X1    g077(.A(new_n265_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n264_), .A2(KEYINPUT68), .A3(new_n265_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT67), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT67), .B1(new_n246_), .B2(new_n248_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n281_), .B(new_n282_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n250_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(KEYINPUT8), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n264_), .A2(new_n265_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n276_), .B(new_n250_), .C1(new_n249_), .C2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT66), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n277_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G29gat), .B(G36gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G43gat), .B(G50gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n260_), .A2(new_n292_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n259_), .B(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n292_), .A2(KEYINPUT71), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n277_), .A2(new_n291_), .A3(new_n288_), .A4(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n298_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT75), .B(KEYINPUT15), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n295_), .B(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n244_), .B(new_n296_), .C1(new_n302_), .C2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n242_), .A2(new_n243_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n306_), .ZN(new_n308_));
  AOI211_X1 g107(.A(new_n238_), .B(new_n239_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT36), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n236_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT37), .B1(new_n309_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n237_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n313_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT37), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n310_), .A2(KEYINPUT78), .A3(new_n237_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .A4(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(KEYINPUT77), .B(KEYINPUT37), .C1(new_n309_), .C2(new_n313_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G183gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT82), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT82), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G183gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n329_), .A3(KEYINPUT25), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(KEYINPUT25), .B2(G183gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(KEYINPUT26), .B(G190gat), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT23), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(G183gat), .A3(G190gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n336_), .A2(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT24), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT83), .B1(new_n343_), .B2(new_n340_), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n343_), .A2(KEYINPUT83), .A3(new_n340_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n334_), .A2(new_n341_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G169gat), .ZN(new_n347_));
  INV_X1    g146(.A(G176gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n342_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n336_), .A2(new_n338_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(G190gat), .B1(new_n327_), .B2(new_n329_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n352_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n327_), .A2(new_n329_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT84), .B(new_n353_), .C1(new_n357_), .C2(G190gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n351_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n346_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT30), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G43gat), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n363_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G227gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT85), .ZN(new_n367_));
  INV_X1    g166(.A(G15gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n364_), .A2(new_n365_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT86), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n374_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT86), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G113gat), .B(G120gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT31), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n375_), .A2(new_n378_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n382_), .ZN(new_n384_));
  OAI211_X1 g183(.A(KEYINPUT86), .B(new_n384_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT19), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT98), .B1(new_n353_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT98), .ZN(new_n392_));
  AOI211_X1 g191(.A(new_n392_), .B(new_n389_), .C1(new_n336_), .C2(new_n338_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n350_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(KEYINPUT25), .B(G183gat), .Z(new_n395_));
  OAI21_X1  g194(.A(new_n341_), .B1(new_n332_), .B2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n343_), .A2(KEYINPUT97), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT97), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n342_), .B2(KEYINPUT24), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n397_), .A2(new_n399_), .A3(new_n340_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n394_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G211gat), .B(G218gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT92), .ZN(new_n404_));
  INV_X1    g203(.A(G197gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n404_), .B1(new_n405_), .B2(G204gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(KEYINPUT21), .A3(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G197gat), .B(G204gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n408_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n410_), .A2(KEYINPUT21), .A3(new_n403_), .A4(new_n406_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n403_), .A2(KEYINPUT21), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n388_), .B1(new_n402_), .B2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n360_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(KEYINPUT20), .A3(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n394_), .B2(new_n401_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n346_), .A2(new_n359_), .A3(new_n413_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT20), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n420_), .A2(KEYINPUT99), .A3(new_n388_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT99), .B1(new_n420_), .B2(new_n388_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n417_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G92gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT18), .B(G64gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n425_), .B(new_n426_), .Z(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n427_), .B(new_n417_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(KEYINPUT100), .A3(new_n430_), .ZN(new_n431_));
  OR3_X1    g230(.A1(new_n423_), .A2(KEYINPUT100), .A3(new_n428_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n381_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G155gat), .B(G162gat), .Z(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT88), .ZN(new_n437_));
  INV_X1    g236(.A(G141gat), .ZN(new_n438_));
  INV_X1    g237(.A(G148gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  OAI22_X1  g239(.A1(new_n440_), .A2(KEYINPUT3), .B1(KEYINPUT89), .B2(KEYINPUT2), .ZN(new_n441_));
  NOR3_X1   g240(.A1(KEYINPUT88), .A2(G141gat), .A3(G148gat), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT3), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G141gat), .A2(G148gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n445_));
  OAI22_X1  g244(.A1(new_n442_), .A2(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n445_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n436_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n444_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT1), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n435_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(G141gat), .B2(G148gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT87), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n434_), .B1(new_n449_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n448_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n441_), .A2(new_n446_), .A3(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n459_), .B(new_n381_), .C1(new_n461_), .C2(new_n436_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(KEYINPUT4), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n459_), .B1(new_n461_), .B2(new_n436_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n467_), .A3(new_n434_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n458_), .A2(new_n464_), .A3(new_n462_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G1gat), .B(G29gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(G85gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT0), .B(G57gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n469_), .A2(new_n470_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT33), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT101), .B1(new_n475_), .B2(KEYINPUT33), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT101), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n469_), .A2(new_n470_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n474_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n478_), .B(new_n479_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n463_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n458_), .A2(new_n465_), .A3(new_n462_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n481_), .A3(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n477_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n433_), .A2(new_n476_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT103), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n489_));
  AOI211_X1 g288(.A(KEYINPUT103), .B(new_n474_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n475_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n427_), .A2(KEYINPUT32), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n417_), .B(new_n493_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT20), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n413_), .A2(KEYINPUT94), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n409_), .A2(new_n411_), .A3(new_n497_), .A4(new_n412_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n499_), .B2(new_n402_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT102), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n416_), .B1(new_n500_), .B2(KEYINPUT102), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n388_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n420_), .A2(new_n388_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n493_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n492_), .A2(new_n494_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n487_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G228gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT91), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n499_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n466_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n515_), .A2(KEYINPUT93), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n466_), .B2(KEYINPUT29), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n513_), .B(new_n514_), .C1(new_n517_), .C2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n415_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n512_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT96), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT96), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n520_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n466_), .A2(KEYINPUT29), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G22gat), .B(G50gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G78gat), .B(G106gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n530_), .B1(new_n466_), .B2(KEYINPUT29), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  AOI211_X1 g335(.A(KEYINPUT95), .B(new_n534_), .C1(new_n532_), .C2(new_n535_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n524_), .B(new_n526_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n536_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n526_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n525_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT104), .B1(new_n510_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT104), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n538_), .A2(new_n542_), .ZN(new_n546_));
  AOI211_X1 g345(.A(new_n545_), .B(new_n546_), .C1(new_n487_), .C2(new_n509_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT27), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n431_), .A2(new_n432_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n388_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n503_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(new_n501_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n428_), .B1(new_n553_), .B2(new_n505_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(KEYINPUT27), .A3(new_n430_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(new_n543_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n491_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n386_), .B1(new_n548_), .B2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n550_), .A2(new_n555_), .A3(new_n543_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT105), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n550_), .A2(new_n555_), .A3(new_n543_), .A4(KEYINPUT105), .ZN(new_n563_));
  AND4_X1   g362(.A1(new_n491_), .A2(new_n562_), .A3(new_n386_), .A4(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n233_), .B(new_n325_), .C1(new_n559_), .C2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n260_), .A2(new_n292_), .A3(new_n208_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n208_), .B1(new_n260_), .B2(new_n292_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT70), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n299_), .A2(new_n301_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n260_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n208_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT12), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n568_), .A2(KEYINPUT12), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n567_), .A2(new_n566_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n570_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G120gat), .B(G148gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n570_), .A2(new_n579_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT73), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n589_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n586_), .B(new_n588_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n220_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n295_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n600_), .B2(new_n304_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n220_), .B(new_n295_), .Z(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G169gat), .B(G197gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n608_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT81), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n565_), .A2(new_n599_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n209_), .A3(new_n492_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT38), .ZN(new_n618_));
  INV_X1    g417(.A(new_n494_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n491_), .A2(new_n619_), .A3(new_n507_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n477_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n432_), .B2(new_n431_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n620_), .B1(new_n622_), .B2(new_n476_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n545_), .B1(new_n623_), .B2(new_n546_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n510_), .A2(KEYINPUT104), .A3(new_n543_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n558_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n386_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n564_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n319_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n615_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n232_), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n491_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n618_), .A2(new_n634_), .ZN(G1324gat));
  NAND3_X1  g434(.A1(new_n616_), .A2(new_n210_), .A3(new_n556_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT106), .ZN(new_n637_));
  INV_X1    g436(.A(new_n556_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G8gat), .B1(new_n633_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT39), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n637_), .A2(KEYINPUT40), .A3(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1325gat));
  NAND3_X1  g444(.A1(new_n616_), .A2(new_n368_), .A3(new_n386_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT107), .ZN(new_n647_));
  OAI21_X1  g446(.A(G15gat), .B1(new_n633_), .B2(new_n627_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT41), .Z(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(new_n649_), .A3(KEYINPUT108), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  OAI21_X1  g453(.A(G22gat), .B1(new_n633_), .B2(new_n543_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT42), .ZN(new_n656_));
  INV_X1    g455(.A(G22gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n616_), .A2(new_n657_), .A3(new_n546_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1327gat));
  INV_X1    g458(.A(new_n233_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n596_), .A2(new_n614_), .A3(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n628_), .A2(new_n629_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G29gat), .B1(new_n662_), .B2(new_n492_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  INV_X1    g463(.A(new_n325_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n664_), .B(new_n665_), .C1(new_n559_), .C2(new_n564_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n628_), .B2(new_n325_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n661_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n632_), .A2(KEYINPUT109), .A3(new_n660_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AND4_X1   g472(.A1(KEYINPUT110), .A2(new_n668_), .A3(KEYINPUT44), .A4(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n672_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT110), .B1(new_n675_), .B2(KEYINPUT44), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n668_), .A2(new_n673_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n680_), .A2(G29gat), .A3(new_n492_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n663_), .B1(new_n677_), .B2(new_n681_), .ZN(G1328gat));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(KEYINPUT111), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n556_), .B(new_n680_), .C1(new_n674_), .C2(new_n676_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G36gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(KEYINPUT111), .ZN(new_n688_));
  NOR4_X1   g487(.A1(new_n628_), .A2(new_n661_), .A3(G36gat), .A4(new_n629_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n556_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n689_), .B2(new_n556_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n685_), .B1(new_n687_), .B2(new_n694_), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n684_), .B(new_n693_), .C1(new_n686_), .C2(G36gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1329gat));
  AOI21_X1  g496(.A(new_n363_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n698_), .B(new_n386_), .C1(new_n674_), .C2(new_n676_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n662_), .A2(new_n386_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n363_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g502(.A(G50gat), .B1(new_n662_), .B2(new_n546_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n677_), .A2(G50gat), .A3(new_n680_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n546_), .ZN(G1331gat));
  NOR2_X1   g505(.A1(new_n598_), .A2(new_n614_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n631_), .A3(new_n233_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n709_), .A2(G57gat), .A3(new_n492_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n596_), .A2(new_n614_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n565_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n492_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n710_), .A2(new_n714_), .ZN(G1332gat));
  INV_X1    g514(.A(new_n713_), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n716_), .A2(G64gat), .A3(new_n638_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n709_), .A2(new_n556_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G64gat), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT112), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n718_), .A2(new_n722_), .A3(G64gat), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n721_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n717_), .B1(new_n724_), .B2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n708_), .B2(new_n627_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n627_), .A2(G71gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n716_), .B2(new_n729_), .ZN(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n708_), .B2(new_n543_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n543_), .A2(G78gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n716_), .B2(new_n733_), .ZN(G1335gat));
  NOR2_X1   g533(.A1(new_n628_), .A2(new_n629_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n707_), .A2(new_n660_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n492_), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n233_), .B(new_n712_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n492_), .A2(G85gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(G1336gat));
  AOI21_X1  g539(.A(G92gat), .B1(new_n736_), .B2(new_n556_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n556_), .A2(G92gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n738_), .B2(new_n742_), .ZN(G1337gat));
  NAND3_X1  g542(.A1(new_n736_), .A2(new_n386_), .A3(new_n254_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT113), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n263_), .B1(new_n738_), .B2(new_n386_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g547(.A1(new_n736_), .A2(new_n256_), .A3(new_n546_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n668_), .A2(new_n546_), .A3(new_n660_), .A4(new_n711_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G106gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G106gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g554(.A(G113gat), .ZN(new_n756_));
  AND4_X1   g555(.A1(new_n492_), .A2(new_n562_), .A3(new_n386_), .A4(new_n563_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n614_), .A2(new_n588_), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n302_), .A2(new_n574_), .B1(KEYINPUT12), .B2(new_n568_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n566_), .B1(new_n760_), .B2(new_n567_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n567_), .A2(new_n566_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n760_), .B2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n576_), .A2(KEYINPUT55), .A3(new_n578_), .A4(new_n577_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n585_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT115), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT56), .B1(new_n766_), .B2(new_n585_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n766_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n759_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n605_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n606_), .A2(new_n603_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n611_), .C1(new_n603_), .C2(new_n602_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n758_), .B(new_n629_), .C1(new_n776_), .C2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n772_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n783_));
  AOI211_X1 g582(.A(KEYINPUT115), .B(KEYINPUT56), .C1(new_n766_), .C2(new_n585_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n775_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n759_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n781_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT57), .B1(new_n787_), .B2(new_n630_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n782_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n780_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n775_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n588_), .B(new_n790_), .C1(new_n791_), .C2(new_n771_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT58), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n665_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n232_), .B1(new_n789_), .B2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n325_), .A2(new_n615_), .A3(new_n596_), .A4(new_n233_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n757_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n797_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n796_), .B(new_n800_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n782_), .A2(new_n788_), .B1(new_n665_), .B2(new_n793_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n233_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT59), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n757_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n799_), .A2(KEYINPUT59), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n756_), .B1(new_n807_), .B2(new_n614_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n799_), .A2(G113gat), .A3(new_n615_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT116), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  INV_X1    g610(.A(new_n809_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n801_), .B1(new_n802_), .B2(new_n232_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n804_), .B1(new_n813_), .B2(new_n757_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n789_), .A2(new_n794_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n660_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n805_), .B1(new_n816_), .B2(new_n801_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n814_), .A2(new_n817_), .A3(new_n615_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n811_), .B(new_n812_), .C1(new_n818_), .C2(new_n756_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n810_), .A2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(new_n807_), .ZN(new_n821_));
  OAI21_X1  g620(.A(G120gat), .B1(new_n821_), .B2(new_n598_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n799_), .ZN(new_n823_));
  INV_X1    g622(.A(G120gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n596_), .B2(KEYINPUT60), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n823_), .B(new_n825_), .C1(KEYINPUT60), .C2(new_n824_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n826_), .A2(KEYINPUT117), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(KEYINPUT117), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n822_), .B1(new_n827_), .B2(new_n828_), .ZN(G1341gat));
  AOI21_X1  g628(.A(G127gat), .B1(new_n823_), .B2(new_n233_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT118), .B(G127gat), .Z(new_n831_));
  NOR2_X1   g630(.A1(new_n821_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n832_), .B2(new_n232_), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n807_), .B2(new_n665_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n799_), .A2(G134gat), .A3(new_n629_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT119), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  INV_X1    g637(.A(new_n836_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n814_), .A2(new_n817_), .A3(new_n325_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n838_), .B(new_n839_), .C1(new_n840_), .C2(new_n834_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n841_), .ZN(G1343gat));
  AND2_X1   g641(.A1(new_n813_), .A2(new_n627_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n843_), .A2(new_n492_), .A3(new_n557_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n438_), .A3(new_n614_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n492_), .A3(new_n557_), .ZN(new_n846_));
  OAI21_X1  g645(.A(G141gat), .B1(new_n846_), .B2(new_n615_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1344gat));
  NAND3_X1  g647(.A1(new_n844_), .A2(new_n439_), .A3(new_n599_), .ZN(new_n849_));
  OAI21_X1  g648(.A(G148gat), .B1(new_n846_), .B2(new_n598_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1345gat));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n844_), .B2(new_n233_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n852_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n846_), .A2(new_n660_), .A3(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1346gat));
  AOI21_X1  g655(.A(G162gat), .B1(new_n844_), .B2(new_n630_), .ZN(new_n857_));
  INV_X1    g656(.A(G162gat), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n846_), .A2(new_n858_), .A3(new_n325_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1347gat));
  NOR2_X1   g659(.A1(new_n638_), .A2(new_n492_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n861_), .A2(new_n386_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n803_), .A2(new_n543_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT122), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n803_), .A2(new_n865_), .A3(new_n543_), .A4(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n614_), .A2(new_n347_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT123), .Z(new_n868_));
  NAND3_X1  g667(.A1(new_n864_), .A2(new_n866_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n862_), .A2(new_n614_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT120), .Z(new_n871_));
  AOI21_X1  g670(.A(new_n233_), .B1(new_n789_), .B2(new_n794_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n543_), .B(new_n871_), .C1(new_n872_), .C2(new_n798_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT121), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n803_), .A2(new_n875_), .A3(new_n543_), .A4(new_n871_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(G169gat), .A3(new_n876_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n877_), .A2(KEYINPUT62), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(KEYINPUT62), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n869_), .B1(new_n878_), .B2(new_n879_), .ZN(G1348gat));
  NAND4_X1  g679(.A1(new_n864_), .A2(new_n594_), .A3(new_n595_), .A4(new_n866_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n813_), .A2(new_n543_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n882_), .A2(G176gat), .A3(new_n599_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n881_), .A2(new_n348_), .B1(new_n883_), .B2(new_n862_), .ZN(G1349gat));
  AND4_X1   g683(.A1(new_n232_), .A2(new_n864_), .A3(new_n395_), .A4(new_n866_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n357_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n882_), .A2(new_n233_), .A3(new_n862_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1350gat));
  NAND3_X1  g687(.A1(new_n864_), .A2(new_n665_), .A3(new_n866_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G190gat), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n864_), .A2(new_n333_), .A3(new_n630_), .A4(new_n866_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1351gat));
  NAND4_X1  g691(.A1(new_n813_), .A2(new_n627_), .A3(new_n546_), .A4(new_n861_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n615_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT124), .B(G197gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1352gat));
  INV_X1    g695(.A(new_n893_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n599_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g698(.A(new_n232_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NOR4_X1   g701(.A1(new_n893_), .A2(new_n900_), .A3(new_n901_), .A4(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n897_), .A2(new_n232_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n901_), .ZN(G1354gat));
  AND3_X1   g704(.A1(new_n813_), .A2(new_n627_), .A3(new_n546_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n630_), .A4(new_n861_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT126), .B(G218gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT125), .B1(new_n893_), .B2(new_n629_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n325_), .A2(new_n909_), .ZN(new_n912_));
  XOR2_X1   g711(.A(new_n912_), .B(KEYINPUT127), .Z(new_n913_));
  NAND2_X1  g712(.A1(new_n897_), .A2(new_n913_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n911_), .A2(new_n914_), .ZN(G1355gat));
endmodule


