//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT6), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G92gat), .Z(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n207_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n216_), .A2(new_n220_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT67), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n216_), .A2(new_n220_), .ZN(new_n225_));
  AND2_X1   g024(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n224_), .B(new_n225_), .C1(new_n228_), .C2(new_n216_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(new_n206_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G85gat), .B(G92gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n215_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n221_), .A2(new_n222_), .ZN(new_n234_));
  AOI211_X1 g033(.A(KEYINPUT8), .B(new_n231_), .C1(new_n234_), .C2(new_n206_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n214_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G36gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G29gat), .ZN(new_n238_));
  INV_X1    g037(.A(G29gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G36gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT73), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n241_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n244_));
  OAI21_X1  g043(.A(G43gat), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n238_), .A2(new_n240_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT73), .ZN(new_n247_));
  INV_X1    g046(.A(G43gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n242_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n245_), .A2(new_n249_), .A3(G50gat), .ZN(new_n250_));
  AOI21_X1  g049(.A(G50gat), .B1(new_n245_), .B2(new_n249_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G50gat), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n243_), .A2(new_n244_), .A3(G43gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n248_), .B1(new_n247_), .B2(new_n242_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n254_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n245_), .A2(new_n249_), .A3(G50gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT15), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n236_), .B1(new_n253_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT34), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT35), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n250_), .A2(new_n251_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n266_), .B(new_n214_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n260_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n257_), .A2(new_n258_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n252_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n257_), .A2(KEYINPUT15), .A3(new_n258_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT74), .B1(new_n272_), .B2(new_n236_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n263_), .A2(new_n264_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n268_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n260_), .A2(KEYINPUT74), .A3(new_n267_), .A4(new_n274_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G190gat), .B(G218gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G134gat), .B(G162gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT36), .Z(new_n281_));
  NAND3_X1  g080(.A1(new_n276_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n280_), .A2(KEYINPUT36), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AOI211_X1 g083(.A(KEYINPUT75), .B(new_n284_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n260_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n275_), .B1(new_n260_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n277_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(new_n290_), .B2(new_n283_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n282_), .B1(new_n285_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT37), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(KEYINPUT76), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n276_), .A2(new_n296_), .A3(new_n277_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n281_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT37), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n298_), .B(new_n299_), .C1(new_n291_), .C2(new_n285_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n293_), .A2(new_n294_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n294_), .B1(new_n293_), .B2(new_n300_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT78), .B(G8gat), .ZN(new_n304_));
  INV_X1    g103(.A(G1gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT14), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G15gat), .B(G22gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G1gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n309_), .A2(G8gat), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(G8gat), .B1(new_n309_), .B2(new_n310_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(G231gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n316_));
  OR2_X1    g115(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G78gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(G78gat), .A3(new_n318_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G57gat), .B(G64gat), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n321_), .B(new_n322_), .C1(KEYINPUT11), .C2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G64gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G57gat), .ZN(new_n326_));
  INV_X1    g125(.A(G57gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G64gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT11), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT69), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n323_), .A2(new_n331_), .A3(KEYINPUT11), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n324_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n324_), .A2(new_n333_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n316_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(KEYINPUT70), .A3(new_n334_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n315_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G127gat), .B(G155gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G183gat), .B(G211gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n315_), .A2(new_n340_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n341_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n338_), .A2(new_n334_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n315_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n315_), .A2(new_n353_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n346_), .B(KEYINPUT17), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n303_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT19), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(KEYINPUT24), .A3(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n365_), .A2(KEYINPUT89), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(KEYINPUT89), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT23), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G183gat), .A3(G190gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n363_), .A2(KEYINPUT24), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n367_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT26), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT88), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n375_), .A2(KEYINPUT26), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT85), .B(G183gat), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n378_), .B(new_n379_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G183gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(KEYINPUT86), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT86), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT25), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n383_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT87), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n366_), .B(new_n374_), .C1(new_n382_), .C2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n381_), .A2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT91), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n372_), .A2(KEYINPUT90), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT90), .B1(new_n368_), .B2(KEYINPUT23), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n391_), .B(new_n392_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT22), .B(G169gat), .ZN(new_n396_));
  INV_X1    g195(.A(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n364_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n394_), .B1(new_n372_), .B2(KEYINPUT90), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT91), .B1(new_n401_), .B2(new_n390_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n395_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G211gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(G218gat), .ZN(new_n405_));
  INV_X1    g204(.A(G218gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(G211gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT21), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT21), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G197gat), .B(G204gat), .Z(new_n412_));
  NAND3_X1  g211(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G197gat), .B(G204gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n414_), .A3(KEYINPUT21), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n389_), .A2(new_n403_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n379_), .A2(new_n376_), .ZN(new_n419_));
  XOR2_X1   g218(.A(KEYINPUT25), .B(G183gat), .Z(new_n420_));
  OAI211_X1 g219(.A(new_n373_), .B(new_n365_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n369_), .A2(new_n371_), .B1(new_n383_), .B2(new_n375_), .ZN(new_n422_));
  OAI22_X1  g221(.A1(new_n421_), .A2(new_n401_), .B1(new_n399_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n413_), .A2(new_n415_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n418_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n362_), .B1(new_n417_), .B2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT20), .B(new_n362_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n389_), .A2(new_n403_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(new_n424_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G8gat), .B(G36gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT18), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(new_n325_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n325_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G92gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n433_), .A3(G92gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OR3_X1    g237(.A1(new_n426_), .A2(new_n429_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT27), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT103), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT20), .B1(new_n423_), .B2(new_n424_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT102), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT102), .B(KEYINPUT20), .C1(new_n423_), .C2(new_n424_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n416_), .B1(new_n389_), .B2(new_n403_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n361_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n417_), .A2(new_n362_), .A3(new_n425_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n442_), .B1(new_n451_), .B2(new_n438_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n439_), .A2(KEYINPUT27), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n451_), .A2(new_n442_), .A3(new_n438_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n441_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G141gat), .B(G148gat), .Z(new_n457_));
  NAND3_X1  g256(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G155gat), .B(G162gat), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n457_), .B(new_n458_), .C1(KEYINPUT1), .C2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT2), .ZN(new_n461_));
  INV_X1    g260(.A(G141gat), .ZN(new_n462_));
  INV_X1    g261(.A(G148gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT3), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G141gat), .A2(G148gat), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n464_), .B(new_n465_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT94), .B1(G141gat), .B2(G148gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n466_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(KEYINPUT94), .A2(G141gat), .A3(G148gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT95), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT94), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT95), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n466_), .A4(new_n469_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n468_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n460_), .B1(new_n477_), .B2(new_n459_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n416_), .B1(new_n478_), .B2(KEYINPUT29), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G228gat), .A2(G233gat), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n480_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G78gat), .B(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT97), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n479_), .A2(new_n480_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n479_), .A2(new_n480_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n483_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT29), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(new_n460_), .C1(new_n477_), .C2(new_n459_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G22gat), .B(G50gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT28), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n481_), .A2(KEYINPUT97), .A3(new_n482_), .A4(new_n484_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n487_), .A2(new_n490_), .A3(new_n497_), .A4(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n490_), .A2(new_n485_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n497_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G127gat), .B(G134gat), .Z(new_n505_));
  XOR2_X1   g304(.A(G113gat), .B(G120gat), .Z(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT31), .Z(new_n508_));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n428_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n389_), .A2(new_n403_), .A3(KEYINPUT30), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G71gat), .B(G99gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G15gat), .B(G43gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n508_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G227gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT92), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT93), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n510_), .A2(new_n511_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n514_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n508_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n516_), .A3(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n519_), .A2(new_n522_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n522_), .B1(new_n519_), .B2(new_n526_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n504_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n498_), .A2(new_n490_), .A3(new_n497_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n531_), .A2(new_n487_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n519_), .A2(new_n526_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n522_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n535_), .A3(new_n527_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G1gat), .B(G29gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT0), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(new_n327_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n210_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT99), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n477_), .A2(new_n459_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT98), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n507_), .A4(new_n460_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n544_), .B(new_n460_), .C1(new_n477_), .C2(new_n459_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n507_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G225gat), .A2(G233gat), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n542_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n550_), .ZN(new_n552_));
  AOI211_X1 g351(.A(KEYINPUT99), .B(new_n552_), .C1(new_n545_), .C2(new_n548_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT4), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n478_), .A2(new_n555_), .A3(new_n507_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n546_), .B(new_n507_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n552_), .B(new_n556_), .C1(new_n557_), .C2(new_n555_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n541_), .B1(new_n554_), .B2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT99), .B1(new_n557_), .B2(new_n552_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n549_), .A2(new_n542_), .A3(new_n550_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n558_), .A2(new_n560_), .A3(new_n541_), .A4(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n456_), .A2(new_n530_), .A3(new_n536_), .A4(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n439_), .A2(new_n440_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n550_), .B(new_n556_), .C1(new_n557_), .C2(new_n555_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT101), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n540_), .B1(new_n557_), .B2(new_n550_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT100), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n549_), .A2(KEYINPUT4), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n573_), .A2(KEYINPUT101), .A3(new_n550_), .A4(new_n556_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n540_), .B(KEYINPUT100), .C1(new_n557_), .C2(new_n550_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n569_), .A2(new_n572_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT33), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n562_), .A2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n554_), .A2(KEYINPUT33), .A3(new_n541_), .A4(new_n558_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n566_), .A2(new_n576_), .A3(new_n578_), .A4(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n436_), .A2(KEYINPUT32), .A3(new_n437_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n581_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n451_), .B2(new_n581_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n559_), .B2(new_n563_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n528_), .A2(new_n529_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n586_), .A3(new_n532_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n565_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n359_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n353_), .B(new_n214_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n337_), .A2(new_n339_), .A3(KEYINPUT12), .ZN(new_n592_));
  INV_X1    g391(.A(new_n236_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G230gat), .ZN(new_n595_));
  INV_X1    g394(.A(G233gat), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n353_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n600_), .B2(new_n236_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n594_), .A2(new_n597_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n593_), .A2(new_n353_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n591_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n597_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(G120gat), .B(G148gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT72), .B(G204gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT5), .B(G176gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n603_), .A2(new_n606_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n590_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n614_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(KEYINPUT13), .A3(new_n612_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n313_), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT81), .B1(new_n620_), .B2(new_n266_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n266_), .B2(new_n620_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n313_), .A2(KEYINPUT81), .A3(new_n269_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n622_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n272_), .A2(new_n313_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n620_), .A2(new_n266_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT82), .B1(new_n629_), .B2(new_n624_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT82), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n627_), .A2(new_n628_), .A3(new_n631_), .A4(new_n623_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G169gat), .B(G197gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT84), .B(G141gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT83), .B(G113gat), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n636_), .B(new_n637_), .Z(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n626_), .A2(new_n630_), .A3(new_n632_), .A4(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n619_), .A2(new_n642_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n589_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n644_), .A2(G1gat), .A3(new_n564_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(KEYINPUT38), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT104), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(KEYINPUT38), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n643_), .A2(new_n358_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n285_), .A2(new_n291_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n298_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n587_), .B2(new_n565_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n654_), .B2(new_n564_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n647_), .A2(new_n648_), .A3(new_n655_), .ZN(G1324gat));
  INV_X1    g455(.A(new_n644_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n456_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n304_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G8gat), .B1(new_n654_), .B2(new_n456_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT39), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT105), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n659_), .A2(new_n661_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(G1325gat));
  OR3_X1    g467(.A1(new_n644_), .A2(G15gat), .A3(new_n586_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G15gat), .B1(new_n654_), .B2(new_n586_), .ZN(new_n673_));
  XOR2_X1   g472(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n672_), .A3(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n654_), .B2(new_n532_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n532_), .A2(G22gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n644_), .B2(new_n679_), .ZN(G1327gat));
  NAND3_X1  g479(.A1(new_n619_), .A2(new_n642_), .A3(new_n358_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n651_), .B1(new_n565_), .B2(new_n587_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n564_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G29gat), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n293_), .A2(new_n300_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT77), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n293_), .A2(new_n294_), .A3(new_n300_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n588_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT43), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n690_), .A2(new_n588_), .A3(new_n694_), .A4(new_n691_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n681_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n688_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  AOI211_X1 g497(.A(KEYINPUT108), .B(new_n681_), .C1(new_n693_), .C2(new_n695_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n687_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n694_), .B1(new_n303_), .B2(new_n588_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n695_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n682_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT108), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n696_), .A2(new_n697_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(KEYINPUT109), .A4(new_n688_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n700_), .A2(new_n706_), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n239_), .B(new_n564_), .C1(new_n696_), .C2(KEYINPUT44), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n686_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  XOR2_X1   g508(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n710_));
  NAND2_X1  g509(.A1(new_n696_), .A2(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n658_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n700_), .B2(new_n706_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n237_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n456_), .A2(G36gat), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n684_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n710_), .B1(new_n714_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  INV_X1    g519(.A(new_n712_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT44), .B1(new_n703_), .B2(KEYINPUT108), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT109), .B1(new_n722_), .B2(new_n705_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n698_), .A2(new_n687_), .A3(new_n699_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G36gat), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n718_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n720_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n720_), .B(new_n728_), .C1(new_n713_), .C2(new_n237_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n719_), .B1(new_n729_), .B2(new_n731_), .ZN(G1329gat));
  INV_X1    g531(.A(new_n586_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G43gat), .B1(new_n684_), .B2(new_n733_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n248_), .B(new_n586_), .C1(new_n696_), .C2(KEYINPUT44), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n707_), .B2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g536(.A1(new_n684_), .A2(new_n254_), .A3(new_n504_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n707_), .A2(new_n504_), .A3(new_n711_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n740_));
  OAI21_X1  g539(.A(G50gat), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n740_), .A2(new_n707_), .A3(new_n504_), .A4(new_n711_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1331gat));
  INV_X1    g542(.A(new_n642_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n618_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n359_), .A2(new_n588_), .A3(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n327_), .B1(new_n747_), .B2(new_n564_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT113), .ZN(new_n749_));
  INV_X1    g548(.A(new_n358_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n653_), .A2(new_n746_), .A3(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT114), .B(G57gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n685_), .A3(new_n752_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n749_), .A2(new_n753_), .ZN(G1332gat));
  AOI21_X1  g553(.A(new_n325_), .B1(new_n751_), .B2(new_n658_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT48), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n658_), .A2(new_n325_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n747_), .B2(new_n757_), .ZN(G1333gat));
  INV_X1    g557(.A(G71gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n751_), .B2(new_n733_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT49), .Z(new_n761_));
  NAND2_X1  g560(.A1(new_n733_), .A2(new_n759_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n747_), .B2(new_n762_), .ZN(G1334gat));
  AOI21_X1  g562(.A(new_n320_), .B1(new_n751_), .B2(new_n504_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT50), .Z(new_n765_));
  NAND2_X1  g564(.A1(new_n504_), .A2(new_n320_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n747_), .B2(new_n766_), .ZN(G1335gat));
  NOR2_X1   g566(.A1(new_n745_), .A2(new_n750_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n683_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n210_), .A3(new_n685_), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n750_), .B(new_n745_), .C1(new_n693_), .C2(new_n695_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(new_n685_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n771_), .B1(new_n773_), .B2(new_n210_), .ZN(G1336gat));
  AOI21_X1  g573(.A(G92gat), .B1(new_n770_), .B2(new_n658_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n456_), .A2(new_n209_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n772_), .B2(new_n776_), .ZN(G1337gat));
  AND2_X1   g576(.A1(new_n772_), .A2(new_n733_), .ZN(new_n778_));
  INV_X1    g577(.A(G99gat), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n733_), .A2(new_n202_), .ZN(new_n780_));
  OAI22_X1  g579(.A1(new_n778_), .A2(new_n779_), .B1(new_n769_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n770_), .A2(new_n203_), .A3(new_n504_), .ZN(new_n783_));
  INV_X1    g582(.A(G106gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n772_), .A2(new_n504_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(KEYINPUT115), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n772_), .A2(new_n788_), .A3(new_n504_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n783_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT53), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n783_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1339gat));
  INV_X1    g595(.A(new_n611_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n597_), .B1(new_n594_), .B2(new_n601_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n602_), .B1(KEYINPUT55), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n594_), .A2(new_n800_), .A3(new_n601_), .A4(new_n597_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT56), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n797_), .C1(new_n799_), .C2(new_n801_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n803_), .A2(new_n642_), .A3(new_n612_), .A4(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n622_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n638_), .C1(new_n623_), .C2(new_n629_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(new_n641_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n651_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n651_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n803_), .A2(new_n809_), .A3(new_n612_), .A4(new_n805_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n613_), .B1(new_n802_), .B2(KEYINPUT56), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n819_), .A2(KEYINPUT58), .A3(new_n809_), .A4(new_n805_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n818_), .A2(new_n690_), .A3(new_n691_), .A4(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n814_), .A2(new_n815_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n358_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n618_), .A2(new_n642_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n750_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT54), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n690_), .A2(new_n691_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n750_), .A4(new_n824_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n823_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n658_), .A2(new_n564_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n733_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n532_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT59), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n504_), .B1(new_n823_), .B2(new_n830_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n834_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n836_), .A2(G113gat), .A3(new_n642_), .A4(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(new_n642_), .A3(new_n834_), .ZN(new_n841_));
  INV_X1    g640(.A(G113gat), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n841_), .A2(KEYINPUT116), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT116), .B1(new_n841_), .B2(new_n842_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n840_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n840_), .B(KEYINPUT117), .C1(new_n843_), .C2(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1340gat));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n838_), .B1(new_n837_), .B2(new_n834_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n822_), .A2(new_n358_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n853_));
  NOR4_X1   g652(.A1(new_n853_), .A2(KEYINPUT59), .A3(new_n504_), .A4(new_n833_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n851_), .B1(new_n855_), .B2(new_n618_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n835_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n619_), .A2(G120gat), .ZN(new_n858_));
  MUX2_X1   g657(.A(new_n858_), .B(G120gat), .S(KEYINPUT60), .Z(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n850_), .B1(new_n856_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n836_), .A2(new_n839_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G120gat), .B1(new_n863_), .B2(new_n619_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(KEYINPUT118), .A3(new_n860_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1341gat));
  AOI21_X1  g665(.A(G127gat), .B1(new_n857_), .B2(new_n750_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n750_), .A2(G127gat), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT119), .Z(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n855_), .B2(new_n869_), .ZN(G1342gat));
  AOI21_X1  g669(.A(G134gat), .B1(new_n857_), .B2(new_n652_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(KEYINPUT120), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(KEYINPUT120), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n303_), .A2(G134gat), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n872_), .A2(new_n873_), .B1(new_n855_), .B2(new_n874_), .ZN(G1343gat));
  NOR3_X1   g674(.A1(new_n853_), .A2(new_n733_), .A3(new_n532_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n832_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n744_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT121), .B(G141gat), .Z(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1344gat));
  NOR2_X1   g679(.A1(new_n877_), .A2(new_n619_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n463_), .ZN(G1345gat));
  NOR2_X1   g681(.A1(new_n877_), .A2(new_n358_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT61), .B(G155gat), .Z(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  OAI21_X1  g684(.A(G162gat), .B1(new_n877_), .B2(new_n827_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n651_), .A2(G162gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n877_), .B2(new_n887_), .ZN(G1347gat));
  NAND2_X1  g687(.A1(new_n831_), .A2(new_n532_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n456_), .A2(new_n685_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n733_), .ZN(new_n891_));
  XOR2_X1   g690(.A(new_n891_), .B(KEYINPUT122), .Z(new_n892_));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n642_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n894_), .A2(G169gat), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n894_), .B2(G169gat), .ZN(new_n897_));
  INV_X1    g696(.A(new_n893_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n642_), .A2(new_n396_), .ZN(new_n899_));
  XOR2_X1   g698(.A(new_n899_), .B(KEYINPUT124), .Z(new_n900_));
  OAI22_X1  g699(.A1(new_n896_), .A2(new_n897_), .B1(new_n898_), .B2(new_n900_), .ZN(G1348gat));
  NAND2_X1  g700(.A1(new_n893_), .A2(new_n618_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g702(.A1(new_n898_), .A2(new_n358_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n381_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n904_), .B2(new_n420_), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n898_), .B2(new_n827_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n651_), .A2(new_n419_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n898_), .B2(new_n908_), .ZN(G1351gat));
  NAND2_X1  g708(.A1(new_n876_), .A2(new_n890_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n642_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n618_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g714(.A(new_n358_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT125), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n911_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n918_), .B(new_n919_), .Z(G1354gat));
  NOR2_X1   g719(.A1(new_n910_), .A2(new_n827_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n652_), .A2(new_n406_), .ZN(new_n922_));
  OAI22_X1  g721(.A1(new_n921_), .A2(new_n406_), .B1(new_n910_), .B2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT126), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925_));
  OAI221_X1 g724(.A(new_n925_), .B1(new_n910_), .B2(new_n922_), .C1(new_n921_), .C2(new_n406_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1355gat));
endmodule


