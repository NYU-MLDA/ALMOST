//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_;
  OAI21_X1  g000(.A(KEYINPUT64), .B1(G85gat), .B2(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203_));
  INV_X1    g002(.A(G85gat), .ZN(new_n204_));
  INV_X1    g003(.A(G92gat), .ZN(new_n205_));
  OAI211_X1 g004(.A(new_n202_), .B(new_n203_), .C1(new_n204_), .C2(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NOR3_X1   g007(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT64), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n206_), .B1(new_n209_), .B2(new_n203_), .ZN(new_n210_));
  AND2_X1   g009(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n211_), .A2(new_n212_), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n210_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n224_), .A2(new_n216_), .A3(new_n217_), .A4(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n207_), .A2(new_n208_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(KEYINPUT8), .A3(new_n227_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n220_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT66), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n234_));
  INV_X1    g033(.A(G57gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(G64gat), .ZN(new_n236_));
  INV_X1    g035(.A(G64gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(G57gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(G57gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(G64gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT11), .ZN(new_n242_));
  XOR2_X1   g041(.A(G71gat), .B(G78gat), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G78gat), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n245_), .A2(KEYINPUT11), .A3(new_n240_), .A4(new_n241_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n244_), .A2(KEYINPUT67), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT67), .B1(new_n244_), .B2(new_n246_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n220_), .A2(new_n230_), .A3(new_n250_), .A4(new_n231_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n233_), .A2(new_n249_), .A3(KEYINPUT12), .A4(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n244_), .A2(new_n246_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n232_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT12), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(G230gat), .A2(G233gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n232_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n253_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n252_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n252_), .A2(new_n260_), .A3(KEYINPUT68), .A4(new_n257_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n253_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n255_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n232_), .A2(KEYINPUT65), .A3(new_n254_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n258_), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G204gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G176gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT69), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n263_), .A2(new_n274_), .A3(new_n264_), .A4(new_n269_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n278_), .A2(new_n279_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n277_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT71), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n284_), .B(new_n277_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT13), .B1(new_n283_), .B2(new_n285_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT13), .ZN(new_n290_));
  INV_X1    g089(.A(new_n285_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n278_), .B(new_n279_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n284_), .B1(new_n292_), .B2(new_n277_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n290_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n285_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT72), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n289_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G15gat), .B(G22gat), .ZN(new_n298_));
  INV_X1    g097(.A(G1gat), .ZN(new_n299_));
  INV_X1    g098(.A(G8gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT14), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G8gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G29gat), .B(G36gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G43gat), .B(G50gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n304_), .B(new_n307_), .Z(new_n308_));
  NAND2_X1  g107(.A1(G229gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n307_), .B(KEYINPUT15), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n304_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n304_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n307_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n315_), .A3(new_n309_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G113gat), .B(G141gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G169gat), .ZN(new_n319_));
  INV_X1    g118(.A(G197gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n322_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n297_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G64gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(new_n205_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G226gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT19), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n333_), .B(KEYINPUT93), .Z(new_n334_));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT77), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(G183gat), .A3(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n335_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n341_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G169gat), .ZN(new_n344_));
  INV_X1    g143(.A(G176gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT24), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347_));
  MUX2_X1   g146(.A(new_n346_), .B(KEYINPUT24), .S(new_n347_), .Z(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT25), .B(G183gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(KEYINPUT75), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT75), .B1(new_n351_), .B2(G183gat), .ZN(new_n352_));
  INV_X1    g151(.A(G190gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT26), .B1(new_n353_), .B2(KEYINPUT76), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n353_), .A2(KEYINPUT26), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n352_), .B(new_n354_), .C1(new_n355_), .C2(KEYINPUT76), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n343_), .B(new_n348_), .C1(new_n350_), .C2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT21), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT90), .B(G204gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(new_n320_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G197gat), .A2(G204gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G211gat), .B(G218gat), .Z(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n320_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n358_), .B1(G197gat), .B2(G204gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n360_), .A2(new_n361_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n363_), .A2(KEYINPUT21), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n362_), .A2(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G169gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT22), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT79), .B(G176gat), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n377_));
  OAI22_X1  g176(.A1(new_n376_), .A2(new_n377_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n336_), .A2(new_n338_), .A3(KEYINPUT23), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(KEYINPUT81), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n380_), .A2(KEYINPUT81), .B1(new_n340_), .B2(new_n342_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n379_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n357_), .B(new_n369_), .C1(new_n378_), .C2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT94), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(KEYINPUT20), .ZN(new_n386_));
  INV_X1    g185(.A(new_n348_), .ZN(new_n387_));
  XOR2_X1   g186(.A(KEYINPUT26), .B(G190gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT95), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n389_), .B2(new_n349_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n381_), .A2(new_n382_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n343_), .B1(G183gat), .B2(G190gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT22), .B(G169gat), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n375_), .A2(new_n394_), .B1(G169gat), .B2(G176gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n369_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n386_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n385_), .B1(new_n384_), .B2(KEYINPUT20), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n334_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT96), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n357_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n405_), .B2(new_n398_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n390_), .A2(new_n391_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n333_), .B1(new_n407_), .B2(new_n369_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n403_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n408_), .A3(new_n403_), .ZN(new_n411_));
  AND4_X1   g210(.A1(new_n331_), .A2(new_n402_), .A3(new_n410_), .A4(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n406_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(new_n409_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n331_), .B1(new_n414_), .B2(new_n402_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT99), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT98), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G113gat), .B(G120gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G127gat), .B(G134gat), .Z(new_n423_));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G127gat), .B(G134gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT83), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n422_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n426_), .B(new_n424_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n422_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT97), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n425_), .A2(new_n427_), .A3(new_n422_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT97), .B1(new_n434_), .B2(new_n428_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT3), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G141gat), .A2(G148gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT2), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n442_));
  INV_X1    g241(.A(G155gat), .ZN(new_n443_));
  INV_X1    g242(.A(G162gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n441_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT1), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n448_), .B(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n447_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n439_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(new_n437_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(KEYINPUT87), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT87), .B1(new_n452_), .B2(new_n454_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n449_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n420_), .B1(new_n436_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n457_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n447_), .A2(new_n448_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n460_), .A2(new_n455_), .B1(new_n441_), .B2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(KEYINPUT98), .A3(new_n435_), .A4(new_n433_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n428_), .B(KEYINPUT84), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n431_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n434_), .A2(KEYINPUT85), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n468_), .A3(new_n458_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n459_), .A2(new_n463_), .A3(KEYINPUT4), .A4(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n428_), .A2(KEYINPUT84), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n428_), .A2(KEYINPUT84), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n471_), .A2(new_n472_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT100), .B(KEYINPUT4), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n458_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n419_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n459_), .A2(new_n463_), .A3(new_n469_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n419_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G29gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT0), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(new_n235_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(new_n204_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n480_), .A2(KEYINPUT33), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n470_), .A2(new_n419_), .A3(new_n475_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n484_), .B1(new_n478_), .B2(new_n419_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT101), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT101), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n487_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n479_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n485_), .B1(new_n495_), .B2(new_n476_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT33), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n416_), .A2(new_n486_), .A3(new_n494_), .A4(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n477_), .A2(new_n484_), .A3(new_n479_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT103), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n496_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n480_), .A2(KEYINPUT103), .A3(new_n485_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n400_), .A2(new_n334_), .A3(new_n401_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n333_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n369_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n397_), .A2(KEYINPUT102), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT102), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n407_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n505_), .B1(new_n512_), .B2(new_n406_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT32), .B(new_n331_), .C1(new_n504_), .C2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n414_), .A2(new_n515_), .A3(new_n402_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n502_), .A2(new_n503_), .A3(new_n514_), .A4(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n499_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G228gat), .ZN(new_n519_));
  INV_X1    g318(.A(G233gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n458_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT89), .B1(new_n458_), .B2(KEYINPUT29), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n398_), .B(new_n522_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n458_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n507_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n521_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT29), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n531_), .B(new_n449_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n526_), .A2(new_n530_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n398_), .A2(new_n522_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n462_), .B2(new_n531_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n539_), .B2(new_n523_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n522_), .B1(new_n507_), .B2(new_n528_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n536_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G78gat), .B(G106gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G22gat), .B(G50gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n535_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n535_), .B2(new_n542_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n464_), .A2(new_n468_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n552_));
  OAI211_X1 g351(.A(G227gat), .B(G233gat), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n464_), .A2(new_n468_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT31), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n473_), .A2(new_n550_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G227gat), .A2(G233gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n405_), .A2(KEYINPUT82), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n561_), .B(new_n357_), .C1(new_n378_), .C2(new_n383_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G15gat), .B(G43gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT30), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n560_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G71gat), .B(G99gat), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n567_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n560_), .A2(new_n562_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n564_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n560_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n569_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n559_), .B1(new_n568_), .B2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n553_), .A2(new_n558_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n567_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n572_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n549_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n584_));
  OAI22_X1  g383(.A1(new_n583_), .A2(new_n584_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n535_), .A2(new_n542_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n545_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n575_), .A2(new_n588_), .A3(new_n579_), .A4(new_n546_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n585_), .A2(new_n589_), .B1(new_n503_), .B2(new_n502_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n414_), .A2(new_n402_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n331_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n414_), .A2(new_n331_), .A3(new_n402_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT27), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n592_), .B1(new_n504_), .B2(new_n513_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n596_), .A2(new_n594_), .A3(KEYINPUT27), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n518_), .A2(new_n582_), .B1(new_n590_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT35), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT34), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n259_), .A2(new_n307_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n233_), .A2(new_n312_), .A3(new_n251_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n603_), .A2(new_n600_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n613_));
  OR3_X1    g412(.A1(new_n608_), .A2(new_n609_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n613_), .B(new_n615_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT16), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(G183gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(G211gat), .ZN(new_n622_));
  INV_X1    g421(.A(G183gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n620_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(G211gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT17), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n622_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n622_), .B2(new_n626_), .ZN(new_n629_));
  AND2_X1   g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n304_), .B(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n631_), .A2(new_n253_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n253_), .ZN(new_n633_));
  NOR4_X1   g432(.A1(new_n628_), .A2(new_n629_), .A3(new_n632_), .A4(new_n633_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n631_), .A2(new_n249_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n631_), .A2(new_n249_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n629_), .A3(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT74), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT74), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n634_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n599_), .A2(new_n618_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n327_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n502_), .A2(new_n503_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n518_), .A2(new_n582_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n590_), .A2(new_n598_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n326_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(KEYINPUT104), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n599_), .B2(new_n326_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n288_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n294_), .A2(KEYINPUT72), .A3(new_n295_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT73), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n614_), .A2(new_n657_), .A3(new_n616_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT37), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n641_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n656_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n644_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n653_), .A2(new_n662_), .A3(new_n299_), .A4(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT105), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(KEYINPUT105), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n645_), .B1(new_n668_), .B2(new_n669_), .ZN(G1324gat));
  INV_X1    g469(.A(new_n598_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n327_), .A2(new_n671_), .A3(new_n642_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(G8gat), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n672_), .B2(G8gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n653_), .A2(new_n662_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n300_), .ZN(new_n677_));
  OAI22_X1  g476(.A1(new_n674_), .A2(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g478(.A(new_n580_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n327_), .A2(new_n680_), .A3(new_n642_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G15gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT107), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n684_), .A3(G15gat), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n686_));
  AND3_X1   g485(.A1(new_n683_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n676_), .A2(G15gat), .A3(new_n580_), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(G1326gat));
  OAI21_X1  g489(.A(G22gat), .B1(new_n643_), .B2(new_n549_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT42), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n549_), .A2(G22gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n676_), .B2(new_n693_), .ZN(G1327gat));
  NOR2_X1   g493(.A1(new_n640_), .A2(new_n617_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n656_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n653_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n663_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n649_), .B(new_n641_), .C1(new_n289_), .C2(new_n296_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n656_), .A2(KEYINPUT109), .A3(new_n649_), .A4(new_n641_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n599_), .B2(new_n659_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n590_), .A2(new_n598_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n581_), .B1(new_n499_), .B2(new_n517_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n705_), .B(new_n660_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n704_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n702_), .A2(KEYINPUT44), .A3(new_n703_), .A4(new_n709_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n710_), .A2(G29gat), .A3(new_n663_), .ZN(new_n711_));
  AOI22_X1  g510(.A1(new_n700_), .A2(new_n701_), .B1(new_n704_), .B2(new_n708_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT44), .B1(new_n712_), .B2(new_n703_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n699_), .B1(new_n711_), .B2(new_n714_), .ZN(G1328gat));
  NAND2_X1  g514(.A1(new_n710_), .A2(new_n671_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G36gat), .B1(new_n716_), .B2(new_n713_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n598_), .A2(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n653_), .A2(new_n696_), .A3(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n717_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT46), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT111), .B(new_n725_), .C1(new_n717_), .C2(new_n721_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1329gat));
  NAND3_X1  g526(.A1(new_n710_), .A2(G43gat), .A3(new_n680_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n697_), .A2(new_n580_), .ZN(new_n729_));
  OAI22_X1  g528(.A1(new_n728_), .A2(new_n713_), .B1(G43gat), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g530(.A1(new_n697_), .A2(G50gat), .A3(new_n549_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n549_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n714_), .A2(new_n733_), .A3(new_n710_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(KEYINPUT112), .A3(G50gat), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT112), .B1(new_n734_), .B2(G50gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n732_), .B1(new_n736_), .B2(new_n737_), .ZN(G1331gat));
  NOR2_X1   g537(.A1(new_n656_), .A2(new_n649_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n642_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n644_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(new_n648_), .A3(new_n661_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n663_), .A2(new_n235_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(G1332gat));
  OR3_X1    g543(.A1(new_n742_), .A2(G64gat), .A3(new_n598_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n739_), .A2(new_n671_), .A3(new_n642_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(G64gat), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n746_), .B2(G64gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n745_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n752_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1333gat));
  OAI21_X1  g554(.A(G71gat), .B1(new_n740_), .B2(new_n580_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT49), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n580_), .A2(G71gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n742_), .B2(new_n758_), .ZN(G1334gat));
  OAI21_X1  g558(.A(G78gat), .B1(new_n740_), .B2(new_n549_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT50), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n742_), .A2(G78gat), .A3(new_n549_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT114), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n765_), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1335gat));
  NAND3_X1  g566(.A1(new_n739_), .A2(new_n648_), .A3(new_n695_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n204_), .A3(new_n663_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n709_), .A2(new_n641_), .A3(new_n739_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n772_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n644_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n770_), .B1(new_n775_), .B2(new_n204_), .ZN(G1336gat));
  NAND3_X1  g575(.A1(new_n769_), .A2(new_n205_), .A3(new_n671_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n598_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n205_), .ZN(G1337gat));
  OR4_X1    g578(.A1(new_n212_), .A2(new_n768_), .A3(new_n211_), .A4(new_n580_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n580_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n222_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT51), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n780_), .B(new_n784_), .C1(new_n781_), .C2(new_n222_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n769_), .A2(new_n223_), .A3(new_n733_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n709_), .A2(new_n733_), .A3(new_n739_), .A4(new_n641_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(G106gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n788_), .B2(G106gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n263_), .A2(new_n794_), .A3(new_n264_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n252_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n252_), .A2(new_n257_), .A3(new_n265_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n796_), .A2(KEYINPUT55), .B1(new_n797_), .B2(new_n258_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n275_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT56), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n800_), .A2(new_n649_), .A3(new_n292_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n321_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(KEYINPUT118), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n313_), .A2(new_n315_), .A3(new_n310_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n802_), .B2(KEYINPUT118), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n324_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n617_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n618_), .A2(new_n809_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n795_), .A2(new_n798_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n276_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n815_), .B(new_n275_), .C1(new_n795_), .C2(new_n798_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n806_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n292_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT119), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT58), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT119), .B(new_n822_), .C1(new_n817_), .C2(new_n819_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n823_), .A3(new_n660_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n810_), .A2(new_n812_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n640_), .A2(new_n326_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n294_), .A2(new_n295_), .A3(new_n659_), .A4(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n830_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n825_), .A2(new_n641_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n671_), .A2(new_n644_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n680_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n833_), .A2(new_n733_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836_), .B2(new_n649_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n824_), .A2(new_n812_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n818_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n800_), .A2(new_n649_), .A3(new_n292_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n841_), .B2(new_n617_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n641_), .B1(new_n838_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n831_), .A2(new_n832_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n835_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n549_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(KEYINPUT59), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n845_), .A2(new_n549_), .A3(new_n846_), .A4(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n649_), .A2(G113gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT121), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n837_), .B1(new_n853_), .B2(new_n855_), .ZN(G1340gat));
  NAND3_X1  g655(.A1(new_n849_), .A2(new_n297_), .A3(new_n852_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G120gat), .ZN(new_n858_));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n656_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(KEYINPUT60), .B2(new_n859_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n847_), .B2(new_n861_), .ZN(G1341gat));
  NOR4_X1   g661(.A1(new_n833_), .A2(new_n733_), .A3(new_n641_), .A4(new_n835_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT122), .B1(new_n863_), .B2(G127gat), .ZN(new_n864_));
  INV_X1    g663(.A(G127gat), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n641_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n848_), .A2(KEYINPUT59), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n852_), .B(new_n866_), .C1(new_n836_), .C2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n869_), .B(new_n865_), .C1(new_n847_), .C2(new_n641_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n864_), .A2(new_n868_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n864_), .A2(new_n868_), .A3(KEYINPUT123), .A4(new_n870_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1342gat));
  INV_X1    g674(.A(G134gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n847_), .B2(new_n617_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n877_), .A2(KEYINPUT124), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n849_), .A2(G134gat), .A3(new_n660_), .A4(new_n852_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(KEYINPUT124), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(G1343gat));
  NOR2_X1   g680(.A1(new_n833_), .A2(new_n585_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n834_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n326_), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n656_), .ZN(new_n886_));
  XOR2_X1   g685(.A(new_n886_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g686(.A1(new_n883_), .A2(new_n641_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT61), .B(G155gat), .Z(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1346gat));
  NOR3_X1   g689(.A1(new_n883_), .A2(new_n444_), .A3(new_n659_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n444_), .B1(new_n883_), .B2(new_n617_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n894_), .B(new_n444_), .C1(new_n883_), .C2(new_n617_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n893_), .B2(new_n895_), .ZN(G1347gat));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n671_), .A2(new_n644_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n580_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n649_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n659_), .B1(new_n820_), .B2(KEYINPUT58), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n841_), .A2(new_n811_), .B1(new_n902_), .B2(new_n823_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n640_), .B1(new_n903_), .B2(new_n810_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n830_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n829_), .B(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n549_), .B(new_n901_), .C1(new_n904_), .C2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n907_), .A2(new_n908_), .A3(G169gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n907_), .B2(G169gat), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n733_), .B(new_n900_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n913_));
  OAI211_X1 g712(.A(KEYINPUT126), .B(new_n911_), .C1(new_n913_), .C2(new_n344_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n394_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n897_), .B1(new_n912_), .B2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT126), .B1(new_n913_), .B2(new_n344_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n907_), .A2(new_n908_), .A3(G169gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n918_), .A2(new_n919_), .A3(KEYINPUT62), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n920_), .A2(KEYINPUT127), .A3(new_n915_), .A4(new_n914_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n921_), .ZN(G1348gat));
  NAND3_X1  g721(.A1(new_n845_), .A2(new_n549_), .A3(new_n899_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n923_), .A2(new_n656_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n345_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n375_), .B2(new_n924_), .ZN(G1349gat));
  NOR2_X1   g725(.A1(new_n923_), .A2(new_n641_), .ZN(new_n927_));
  MUX2_X1   g726(.A(G183gat), .B(new_n349_), .S(new_n927_), .Z(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n923_), .B2(new_n659_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n618_), .A2(new_n389_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n923_), .B2(new_n930_), .ZN(G1351gat));
  NAND3_X1  g730(.A1(new_n882_), .A2(new_n644_), .A3(new_n671_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n326_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n320_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n656_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(G204gat), .ZN(new_n936_));
  INV_X1    g735(.A(new_n359_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n935_), .ZN(G1353gat));
  NOR2_X1   g737(.A1(new_n932_), .A2(new_n641_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n939_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(KEYINPUT63), .B(G211gat), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n932_), .A2(new_n641_), .A3(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n940_), .A2(new_n942_), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n932_), .B2(new_n659_), .ZN(new_n944_));
  OR2_X1    g743(.A1(new_n617_), .A2(G218gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n932_), .B2(new_n945_), .ZN(G1355gat));
endmodule


