//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT15), .Z(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G229gat), .A2(G233gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n212_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n204_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n212_), .B(new_n204_), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n213_), .A2(new_n218_), .B1(new_n219_), .B2(new_n215_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G113gat), .B(G141gat), .Z(new_n221_));
  XNOR2_X1  g020(.A(G169gat), .B(G197gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n220_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT12), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT6), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT6), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G99gat), .A3(G106gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n228_), .A2(new_n230_), .A3(KEYINPUT65), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT65), .B1(new_n228_), .B2(new_n230_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  INV_X1    g033(.A(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT9), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(G85gat), .A3(G92gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G85gat), .B(G92gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n237_), .B(new_n239_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n233_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n228_), .A2(new_n230_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246_));
  INV_X1    g045(.A(G99gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n235_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n244_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT8), .B1(new_n251_), .B2(new_n240_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n248_), .A2(new_n249_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n240_), .A2(KEYINPUT8), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n242_), .B1(new_n252_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G71gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(KEYINPUT67), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(KEYINPUT67), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G78gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(G78gat), .B1(new_n259_), .B2(new_n260_), .ZN(new_n264_));
  INV_X1    g063(.A(G64gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G57gat), .ZN(new_n266_));
  INV_X1    g065(.A(G57gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G64gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n268_), .A3(KEYINPUT11), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT11), .B1(new_n266_), .B2(new_n268_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n263_), .B(new_n264_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n264_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n259_), .A2(new_n260_), .A3(G78gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n269_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n226_), .B1(new_n257_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G230gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT64), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n257_), .B2(new_n276_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT8), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n229_), .B1(G99gat), .B2(G106gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n227_), .A2(KEYINPUT6), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT66), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n228_), .A2(new_n230_), .A3(new_n243_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(new_n253_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n240_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n282_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n255_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n228_), .A2(new_n230_), .A3(KEYINPUT65), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n290_), .B1(new_n294_), .B2(new_n253_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n281_), .B1(new_n289_), .B2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n245_), .A2(new_n250_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n240_), .B1(new_n297_), .B2(new_n286_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n256_), .B(KEYINPUT68), .C1(new_n298_), .C2(new_n282_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n242_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n276_), .A2(new_n226_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n277_), .B(new_n280_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n242_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n276_), .B(new_n304_), .C1(new_n289_), .C2(new_n295_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n257_), .A2(new_n276_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n279_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G120gat), .B(G148gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT5), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G176gat), .B(G204gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n303_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT69), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n303_), .A2(new_n308_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n312_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n318_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT71), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n320_), .B(new_n326_), .C1(new_n318_), .C2(new_n323_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n225_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT88), .B(G204gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n330_), .B2(G197gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(G211gat), .B(G218gat), .Z(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(KEYINPUT21), .A3(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT89), .ZN(new_n334_));
  INV_X1    g133(.A(G197gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(G204gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT87), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n330_), .A2(new_n335_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT21), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n332_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n339_), .B(new_n340_), .C1(KEYINPUT21), .C2(new_n331_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT23), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(G183gat), .B2(G190gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G169gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G169gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n350_), .B2(KEYINPUT22), .ZN(new_n351_));
  INV_X1    g150(.A(G176gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n345_), .B(new_n346_), .C1(new_n349_), .C2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n352_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n356_));
  INV_X1    g155(.A(G190gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT26), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT26), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(KEYINPUT76), .A3(G190gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT25), .B(G183gat), .Z(new_n362_));
  INV_X1    g161(.A(KEYINPUT24), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n355_), .A2(new_n346_), .ZN(new_n364_));
  OAI22_X1  g163(.A1(new_n361_), .A2(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n366_));
  OAI221_X1 g165(.A(new_n344_), .B1(KEYINPUT24), .B2(new_n355_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n365_), .A2(new_n366_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n354_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT79), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n371_), .B(new_n354_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n342_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT19), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n334_), .A2(new_n341_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT92), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n345_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n347_), .A2(new_n352_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n346_), .A3(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n345_), .A2(new_n377_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n382_));
  INV_X1    g181(.A(new_n355_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n344_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT26), .B(G190gat), .Z(new_n386_));
  OAI22_X1  g185(.A1(new_n362_), .A2(new_n386_), .B1(new_n364_), .B2(new_n382_), .ZN(new_n387_));
  OAI22_X1  g186(.A1(new_n380_), .A2(new_n381_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT20), .B1(new_n376_), .B2(new_n388_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n373_), .A2(new_n375_), .A3(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n375_), .B(KEYINPUT90), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n370_), .A2(new_n342_), .A3(new_n372_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n376_), .B2(new_n388_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n392_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G8gat), .B(G36gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT18), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT96), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT97), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(KEYINPUT97), .A3(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G155gat), .B(G162gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT2), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT3), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n410_), .B1(new_n419_), .B2(KEYINPUT86), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(KEYINPUT86), .B2(new_n419_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n413_), .B(KEYINPUT84), .ZN(new_n422_));
  AND2_X1   g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n423_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n422_), .B(new_n424_), .C1(KEYINPUT1), .C2(new_n410_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G127gat), .B(G134gat), .Z(new_n427_));
  XOR2_X1   g226(.A(G113gat), .B(G120gat), .Z(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n421_), .A2(new_n425_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n429_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n431_), .B(KEYINPUT4), .C1(KEYINPUT93), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n432_), .A2(new_n435_), .A3(new_n436_), .A4(new_n429_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n409_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n431_), .A2(new_n433_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n409_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G1gat), .B(G29gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(G85gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT0), .B(G57gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  OR3_X1    g244(.A1(new_n438_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n375_), .B1(new_n373_), .B2(new_n389_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n393_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n402_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT98), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n452_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n408_), .A2(new_n448_), .A3(new_n453_), .A4(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT95), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n409_), .B1(new_n439_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n456_), .B2(new_n439_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n445_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n434_), .A2(new_n437_), .A3(new_n409_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n397_), .A2(new_n401_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n401_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(new_n390_), .B2(new_n396_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n447_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT94), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n447_), .A2(new_n466_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n447_), .A2(new_n470_), .A3(new_n466_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n465_), .A2(new_n468_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n455_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G227gat), .A2(G233gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n474_), .B(KEYINPUT80), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT30), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT83), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n479_));
  XOR2_X1   g278(.A(new_n429_), .B(new_n479_), .Z(new_n480_));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT81), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G15gat), .B(G43gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n370_), .A2(new_n372_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n480_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n485_), .A2(new_n486_), .A3(new_n480_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n478_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n489_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(new_n477_), .A3(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n432_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT29), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n376_), .B1(new_n426_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT28), .B1(new_n432_), .B2(KEYINPUT29), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G228gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(new_n262_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(new_n235_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G22gat), .B(G50gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  OR3_X1    g306(.A1(new_n500_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n495_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n473_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n490_), .A2(new_n493_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n448_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n462_), .A2(KEYINPUT27), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n449_), .A2(new_n450_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n463_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n462_), .A2(new_n464_), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT99), .B(KEYINPUT27), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n516_), .A2(new_n518_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n512_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n328_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G190gat), .B(G218gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G134gat), .B(G162gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(KEYINPUT34), .Z(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n531_));
  NOR3_X1   g330(.A1(new_n530_), .A2(KEYINPUT74), .A3(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n530_), .A2(new_n531_), .ZN(new_n533_));
  AOI211_X1 g332(.A(new_n532_), .B(new_n533_), .C1(new_n257_), .C2(new_n217_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n205_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(new_n300_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n530_), .A2(new_n531_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(KEYINPUT74), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT74), .ZN(new_n540_));
  OAI221_X1 g339(.A(new_n534_), .B1(new_n540_), .B2(new_n537_), .C1(new_n535_), .C2(new_n300_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT73), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n528_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n544_), .A2(new_n545_), .B1(new_n528_), .B2(new_n542_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT73), .B1(new_n539_), .B2(new_n541_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT36), .B1(new_n547_), .B2(new_n528_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n546_), .A2(KEYINPUT37), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT37), .B1(new_n546_), .B2(new_n548_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n212_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n272_), .A2(new_n275_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT75), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G127gat), .B(G155gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT16), .ZN(new_n558_));
  XOR2_X1   g357(.A(G183gat), .B(G211gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT17), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n556_), .B(new_n562_), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n555_), .A2(KEYINPUT17), .A3(new_n561_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n551_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n525_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(new_n207_), .A3(new_n448_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT38), .ZN(new_n569_));
  INV_X1    g368(.A(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n328_), .A2(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n571_), .A2(KEYINPUT100), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(KEYINPUT100), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n473_), .A2(new_n511_), .B1(new_n515_), .B2(new_n522_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n546_), .A2(new_n548_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n572_), .A2(new_n573_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n448_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G1gat), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n569_), .A2(new_n580_), .ZN(G1324gat));
  INV_X1    g380(.A(new_n522_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n567_), .A2(new_n208_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT39), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n582_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n585_), .B2(G8gat), .ZN(new_n586_));
  AOI211_X1 g385(.A(KEYINPUT39), .B(new_n208_), .C1(new_n577_), .C2(new_n582_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n583_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT40), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(G1325gat));
  INV_X1    g389(.A(G15gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n567_), .A2(new_n591_), .A3(new_n495_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n495_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G15gat), .B1(new_n578_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT41), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n592_), .B1(new_n596_), .B2(new_n597_), .ZN(G1326gat));
  INV_X1    g397(.A(G22gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n567_), .A2(new_n599_), .A3(new_n510_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n510_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G22gat), .B1(new_n578_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n602_), .A2(new_n603_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n600_), .B1(new_n604_), .B2(new_n605_), .ZN(G1327gat));
  INV_X1    g405(.A(new_n575_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(new_n570_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n525_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(G29gat), .B1(new_n609_), .B2(new_n448_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n524_), .A2(KEYINPUT43), .A3(new_n551_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n575_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n546_), .A2(KEYINPUT37), .A3(new_n548_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n613_), .B1(new_n574_), .B2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(new_n618_), .A3(new_n565_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n325_), .A2(new_n327_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n224_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n611_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n593_), .A2(new_n601_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n472_), .B2(new_n455_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n515_), .A2(new_n522_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n551_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n570_), .B1(new_n626_), .B2(new_n613_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n627_), .A2(KEYINPUT44), .A3(new_n328_), .A4(new_n612_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n622_), .A2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n448_), .A2(G29gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n610_), .B1(new_n629_), .B2(new_n630_), .ZN(G1328gat));
  INV_X1    g430(.A(G36gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n609_), .A2(new_n632_), .A3(new_n582_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT45), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n622_), .A2(new_n628_), .A3(new_n582_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(G36gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT102), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1329gat));
  INV_X1    g438(.A(G43gat), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n593_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n622_), .A2(new_n628_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT103), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n622_), .A2(new_n628_), .A3(new_n644_), .A4(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n328_), .A2(new_n524_), .A3(new_n495_), .A4(new_n608_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n640_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n646_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT106), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n646_), .A2(new_n654_), .A3(new_n651_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n653_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n656_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n646_), .B2(new_n651_), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT106), .B(new_n650_), .C1(new_n643_), .C2(new_n645_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n661_), .ZN(G1330gat));
  AOI21_X1  g461(.A(G50gat), .B1(new_n609_), .B2(new_n510_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n510_), .A2(G50gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n629_), .B2(new_n664_), .ZN(G1331gat));
  INV_X1    g464(.A(new_n620_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n565_), .A2(new_n224_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n576_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n668_), .A2(new_n267_), .A3(new_n579_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT108), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n666_), .A2(new_n225_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n574_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n566_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n579_), .B1(new_n673_), .B2(KEYINPUT107), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(KEYINPUT107), .B2(new_n673_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n670_), .B1(new_n675_), .B2(new_n267_), .ZN(G1332gat));
  OAI21_X1  g475(.A(G64gat), .B1(new_n668_), .B2(new_n522_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT48), .ZN(new_n678_));
  INV_X1    g477(.A(new_n673_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(new_n265_), .A3(new_n582_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1333gat));
  OAI21_X1  g480(.A(G71gat), .B1(new_n668_), .B2(new_n593_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT49), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n679_), .A2(new_n258_), .A3(new_n495_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1334gat));
  OAI21_X1  g484(.A(G78gat), .B1(new_n668_), .B2(new_n601_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT50), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n679_), .A2(new_n262_), .A3(new_n510_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1335gat));
  AND2_X1   g488(.A1(new_n672_), .A2(new_n608_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G85gat), .B1(new_n690_), .B2(new_n448_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT109), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n619_), .A2(new_n671_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT110), .ZN(new_n694_));
  OR3_X1    g493(.A1(new_n619_), .A2(new_n671_), .A3(KEYINPUT110), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n448_), .A2(G85gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n692_), .B1(new_n696_), .B2(new_n697_), .ZN(G1336gat));
  AOI21_X1  g497(.A(G92gat), .B1(new_n690_), .B2(new_n582_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT111), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n696_), .A2(G92gat), .A3(new_n582_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1337gat));
  NAND4_X1  g501(.A1(new_n690_), .A2(new_n234_), .A3(new_n236_), .A4(new_n495_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n593_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n247_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(G1338gat));
  NAND3_X1  g506(.A1(new_n690_), .A2(new_n235_), .A3(new_n510_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n693_), .A2(new_n601_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G106gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G106gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n708_), .B(new_n714_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1339gat));
  NAND2_X1  g517(.A1(new_n315_), .A2(new_n224_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n277_), .B(new_n305_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n303_), .A2(KEYINPUT55), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n296_), .A2(new_n299_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n304_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n301_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT55), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n277_), .A4(new_n280_), .ZN(new_n726_));
  AOI221_X4 g525(.A(KEYINPUT115), .B1(new_n279_), .B2(new_n720_), .C1(new_n721_), .C2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT115), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n721_), .A2(new_n726_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n720_), .A2(new_n279_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n312_), .B1(new_n727_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT56), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(KEYINPUT56), .B(new_n312_), .C1(new_n727_), .C2(new_n731_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n719_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n315_), .A2(new_n317_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n213_), .B(new_n215_), .C1(new_n204_), .C2(new_n212_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n223_), .B1(new_n219_), .B2(new_n214_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n738_), .A2(new_n739_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n737_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n607_), .B1(new_n736_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(KEYINPUT116), .A3(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT58), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n734_), .A2(new_n735_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n315_), .A2(new_n740_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n745_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT58), .B(new_n747_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n551_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT57), .B(new_n607_), .C1(new_n736_), .C2(new_n741_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n744_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT116), .B1(new_n742_), .B2(new_n743_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n565_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n667_), .B(KEYINPUT114), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n617_), .A2(new_n324_), .A3(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT54), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n582_), .A2(new_n579_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n514_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n759_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT59), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n757_), .B(KEYINPUT54), .Z(new_n766_));
  AND2_X1   g565(.A1(new_n742_), .A2(new_n743_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n304_), .B1(new_n289_), .B2(new_n295_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT12), .B1(new_n768_), .B2(new_n554_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n723_), .B2(new_n301_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n725_), .B1(new_n770_), .B2(new_n280_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n303_), .A2(KEYINPUT55), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n730_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT115), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n729_), .A2(new_n728_), .A3(new_n730_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n312_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n735_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n748_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT58), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n746_), .A2(new_n745_), .A3(new_n748_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n617_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT117), .B1(new_n767_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n742_), .A2(new_n743_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT117), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n751_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n752_), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n766_), .B1(new_n787_), .B2(new_n565_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n762_), .A2(KEYINPUT59), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n765_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G113gat), .B1(new_n791_), .B2(new_n225_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n225_), .A2(G113gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n764_), .B2(new_n793_), .ZN(G1340gat));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n791_), .B2(new_n620_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n788_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n789_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n798_), .A2(KEYINPUT118), .A3(new_n666_), .A4(new_n765_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n799_), .A3(G120gat), .ZN(new_n800_));
  INV_X1    g599(.A(new_n764_), .ZN(new_n801_));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n620_), .B2(KEYINPUT60), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n801_), .B(new_n803_), .C1(KEYINPUT60), .C2(new_n802_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n804_), .ZN(G1341gat));
  INV_X1    g604(.A(G127gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n764_), .B2(new_n565_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT119), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n791_), .A2(new_n806_), .A3(new_n565_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1342gat));
  OAI21_X1  g609(.A(G134gat), .B1(new_n791_), .B2(new_n617_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n607_), .A2(G134gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n764_), .B2(new_n812_), .ZN(G1343gat));
  AND2_X1   g612(.A1(new_n755_), .A2(new_n758_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n513_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n760_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n224_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n666_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g620(.A1(new_n816_), .A2(new_n565_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT61), .B(G155gat), .Z(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1346gat));
  OR3_X1    g623(.A1(new_n816_), .A2(G162gat), .A3(new_n607_), .ZN(new_n825_));
  OAI21_X1  g624(.A(G162gat), .B1(new_n816_), .B2(new_n617_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1347gat));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n522_), .A2(new_n448_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n514_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n224_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT120), .B1(new_n788_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834_));
  INV_X1    g633(.A(new_n832_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n752_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n751_), .A2(new_n784_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(KEYINPUT117), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n570_), .B1(new_n838_), .B2(new_n786_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n834_), .B(new_n835_), .C1(new_n839_), .C2(new_n766_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n833_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n797_), .A2(new_n347_), .A3(new_n835_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n835_), .B1(new_n839_), .B2(new_n766_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n350_), .B1(new_n844_), .B2(KEYINPUT120), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT62), .B1(new_n845_), .B2(new_n840_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n828_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n833_), .A2(G169gat), .A3(new_n840_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(KEYINPUT121), .A3(new_n842_), .A4(new_n841_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n851_), .ZN(G1348gat));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n814_), .B2(new_n510_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n759_), .A2(KEYINPUT123), .A3(new_n601_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n830_), .A2(new_n593_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n857_), .A2(new_n352_), .A3(new_n620_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n797_), .A2(new_n831_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n352_), .B1(new_n859_), .B2(new_n620_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT122), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n862_), .B(new_n352_), .C1(new_n859_), .C2(new_n620_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n858_), .B1(new_n861_), .B2(new_n863_), .ZN(G1349gat));
  INV_X1    g663(.A(new_n859_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n865_), .A2(new_n570_), .A3(new_n362_), .ZN(new_n866_));
  AND4_X1   g665(.A1(new_n570_), .A2(new_n854_), .A3(new_n855_), .A4(new_n856_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868_));
  AOI21_X1  g667(.A(G183gat), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT124), .B1(new_n857_), .B2(new_n565_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n866_), .B1(new_n869_), .B2(new_n870_), .ZN(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n859_), .B2(new_n617_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n607_), .A2(new_n386_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n859_), .B2(new_n873_), .ZN(G1351gat));
  NOR3_X1   g673(.A1(new_n814_), .A2(new_n513_), .A3(new_n830_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n224_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n666_), .ZN(new_n878_));
  INV_X1    g677(.A(G204gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n875_), .A2(new_n666_), .A3(new_n330_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1353gat));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n886_));
  INV_X1    g685(.A(G211gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n570_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT126), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n875_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n887_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1354gat));
  AOI21_X1  g691(.A(G218gat), .B1(new_n875_), .B2(new_n575_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n551_), .A2(G218gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT127), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n875_), .B2(new_n895_), .ZN(G1355gat));
endmodule


