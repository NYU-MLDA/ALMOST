//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n212_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n212_), .B(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n217_), .B(new_n213_), .C1(new_n221_), .C2(new_n209_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n219_), .A2(new_n222_), .A3(KEYINPUT74), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT74), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n216_), .A2(new_n224_), .A3(new_n218_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G141gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G197gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n227_), .B(new_n228_), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n229_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n223_), .A2(new_n225_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G176gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n243_));
  INV_X1    g042(.A(G169gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT22), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n244_), .A2(KEYINPUT22), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n242_), .B(new_n245_), .C1(new_n246_), .C2(new_n243_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT24), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n240_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT26), .B(G190gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT25), .B(G183gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n234_), .B(KEYINPUT23), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n241_), .A2(new_n247_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G15gat), .B(G43gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT77), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n258_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT31), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263_));
  INV_X1    g062(.A(G71gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G99gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT76), .B(KEYINPUT30), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269_));
  INV_X1    g068(.A(G120gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(G113gat), .ZN(new_n271_));
  INV_X1    g070(.A(G113gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(G120gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n273_), .A3(KEYINPUT78), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT78), .B1(new_n271_), .B2(new_n273_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n269_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(new_n273_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT78), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n269_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n274_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT79), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n283_), .B2(new_n277_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n268_), .B(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n262_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n262_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT80), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(G155gat), .A3(G162gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT81), .B1(new_n295_), .B2(KEYINPUT1), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n295_), .B2(KEYINPUT1), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n292_), .A2(new_n294_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n296_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT82), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n303_), .A2(KEYINPUT2), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311_));
  AOI22_X1  g110(.A1(KEYINPUT2), .A2(new_n303_), .B1(new_n304_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n295_), .B1(G155gat), .B2(G162gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT83), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n295_), .B(new_n316_), .C1(G155gat), .C2(G162gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n306_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT21), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT88), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT85), .ZN(new_n326_));
  INV_X1    g125(.A(G197gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(G204gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(G204gat), .ZN(new_n329_));
  INV_X1    g128(.A(G204gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n324_), .A2(new_n325_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n325_), .B1(new_n324_), .B2(new_n332_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n322_), .B1(new_n337_), .B2(new_n323_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n328_), .A2(new_n331_), .A3(new_n323_), .A4(new_n329_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n340_), .A2(KEYINPUT86), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(KEYINPUT86), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n339_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT87), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n331_), .A2(new_n329_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT86), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n323_), .A4(new_n328_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n340_), .A2(KEYINPUT86), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n339_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n336_), .B1(new_n344_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G233gat), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n353_), .A2(KEYINPUT84), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(KEYINPUT84), .ZN(new_n355_));
  OAI21_X1  g154(.A(G228gat), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n321_), .A2(new_n352_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n321_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n352_), .A2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n334_), .A2(new_n335_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n350_), .B1(new_n349_), .B2(new_n339_), .ZN(new_n364_));
  AOI211_X1 g163(.A(KEYINPUT87), .B(new_n338_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n363_), .B(new_n361_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n360_), .B1(new_n362_), .B2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT90), .B1(new_n368_), .B2(new_n357_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT89), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n321_), .B1(new_n371_), .B2(new_n366_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT90), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n356_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n359_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT92), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G78gat), .B(G106gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n319_), .A2(new_n320_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n379_), .B(KEYINPUT28), .ZN(new_n384_));
  INV_X1    g183(.A(new_n382_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n368_), .A2(KEYINPUT90), .A3(new_n357_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n373_), .B1(new_n372_), .B2(new_n356_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n358_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n377_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n387_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n378_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT92), .B1(new_n390_), .B2(new_n391_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n389_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n395_), .A2(KEYINPUT91), .A3(new_n391_), .A4(new_n359_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n387_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n375_), .A2(new_n377_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n390_), .A2(new_n391_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n393_), .A2(new_n394_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT18), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n405_), .B(new_n406_), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT32), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n256_), .A2(KEYINPUT94), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n254_), .A2(new_n411_), .A3(new_n255_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n252_), .B(KEYINPUT93), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n250_), .B1(new_n414_), .B2(new_n251_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT22), .B(G169gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n242_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n239_), .A2(KEYINPUT95), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n239_), .A2(KEYINPUT95), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n420_), .A2(KEYINPUT96), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n238_), .B1(new_n420_), .B2(KEYINPUT96), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n413_), .A2(new_n415_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n371_), .A2(new_n366_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT20), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT101), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n258_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n370_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT19), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n352_), .A2(new_n258_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n415_), .A2(new_n413_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n421_), .A2(new_n422_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n370_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n439_), .A3(KEYINPUT20), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n433_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n409_), .B1(new_n434_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G29gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(G85gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT0), .B(G57gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n306_), .A2(new_n318_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n285_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n277_), .A2(new_n282_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT99), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT99), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n277_), .A2(new_n282_), .A3(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n452_), .A2(new_n306_), .A3(new_n318_), .A4(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n449_), .A2(new_n450_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT100), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n450_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT4), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n449_), .B2(new_n455_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT4), .B1(new_n448_), .B2(new_n285_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n459_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n447_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n458_), .A2(new_n447_), .A3(new_n463_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT97), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(new_n370_), .B2(new_n438_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n370_), .B2(new_n428_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n352_), .A2(KEYINPUT97), .A3(new_n423_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n433_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n435_), .A2(new_n439_), .A3(KEYINPUT20), .A4(new_n433_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n465_), .A2(new_n466_), .B1(new_n476_), .B2(new_n408_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n407_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT98), .ZN(new_n479_));
  INV_X1    g278(.A(new_n407_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n475_), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n474_), .A2(KEYINPUT98), .A3(new_n475_), .A4(new_n480_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n450_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n449_), .A2(new_n459_), .A3(new_n455_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n486_), .A2(new_n446_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT33), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n466_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n466_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n442_), .A2(new_n477_), .B1(new_n484_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n290_), .B1(new_n403_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT27), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n482_), .A2(new_n496_), .A3(new_n483_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n465_), .A2(new_n466_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n441_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(new_n407_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT102), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n476_), .B2(new_n407_), .ZN(new_n503_));
  AOI211_X1 g302(.A(KEYINPUT102), .B(new_n480_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT27), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n497_), .B(new_n499_), .C1(new_n501_), .C2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n394_), .A2(new_n378_), .A3(new_n392_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n400_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n508_));
  AOI211_X1 g307(.A(new_n377_), .B(new_n358_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n507_), .B1(new_n510_), .B2(new_n397_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n497_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n498_), .A2(new_n289_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n495_), .A2(new_n512_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT10), .B(G99gat), .Z(new_n517_));
  INV_X1    g316(.A(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G85gat), .B(G92gat), .Z(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT9), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(G85gat), .A3(G92gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT6), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .A4(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT7), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n524_), .B(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n520_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT8), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G85gat), .B(G92gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n527_), .B(KEYINPUT7), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(new_n525_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n212_), .B(new_n526_), .C1(new_n533_), .C2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT34), .Z(new_n541_));
  INV_X1    g340(.A(KEYINPUT35), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n541_), .A2(new_n542_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  AND4_X1   g345(.A1(new_n523_), .A2(new_n519_), .A3(new_n521_), .A4(new_n525_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n532_), .A2(KEYINPUT8), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n536_), .A2(new_n537_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT68), .B1(new_n550_), .B2(new_n221_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n526_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n212_), .B(KEYINPUT15), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n546_), .A2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G190gat), .B(G218gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n559_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT36), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT71), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n544_), .A2(KEYINPUT69), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n539_), .A2(new_n565_), .A3(new_n543_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n556_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n567_), .A2(KEYINPUT70), .A3(new_n545_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT70), .B1(new_n567_), .B2(new_n545_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n557_), .B(new_n563_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT72), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n567_), .A2(new_n545_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n567_), .A2(KEYINPUT70), .A3(new_n545_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n577_), .A2(KEYINPUT72), .A3(new_n557_), .A4(new_n563_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n572_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n557_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n560_), .A2(KEYINPUT36), .A3(new_n561_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n562_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n516_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT64), .B(G71gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(G78gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G57gat), .B(G64gat), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n589_), .A2(KEYINPUT11), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(KEYINPUT11), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n588_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n590_), .B2(new_n588_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n552_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n586_), .B1(new_n594_), .B2(KEYINPUT65), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n552_), .A2(new_n593_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT65), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n552_), .A2(new_n593_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(KEYINPUT12), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n552_), .B2(new_n593_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT66), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n586_), .B1(new_n552_), .B2(new_n593_), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n601_), .A2(new_n603_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n604_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n600_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT5), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n600_), .B(new_n615_), .C1(new_n606_), .C2(new_n608_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(KEYINPUT67), .B(KEYINPUT13), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT13), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n614_), .B(new_n616_), .C1(KEYINPUT67), .C2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n208_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(new_n593_), .Z(new_n625_));
  XOR2_X1   g424(.A(G127gat), .B(G155gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(KEYINPUT17), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n625_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n630_), .B(KEYINPUT17), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n625_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  AND4_X1   g434(.A1(new_n233_), .A2(new_n585_), .A3(new_n622_), .A4(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(new_n498_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n203_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  INV_X1    g438(.A(new_n233_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n579_), .A2(KEYINPUT37), .A3(new_n583_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT37), .B1(new_n579_), .B2(new_n583_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n622_), .A3(new_n635_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n516_), .A2(new_n640_), .A3(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n498_), .A2(KEYINPUT103), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n498_), .A2(KEYINPUT103), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n203_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n638_), .B1(new_n639_), .B2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n650_), .B1(new_n639_), .B2(new_n649_), .ZN(G1324gat));
  NAND3_X1  g450(.A1(new_n645_), .A2(new_n204_), .A3(new_n513_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n636_), .A2(new_n513_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(G8gat), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n653_), .B2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT40), .B(new_n652_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1325gat));
  INV_X1    g460(.A(G15gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n636_), .B2(new_n290_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n645_), .A2(new_n662_), .A3(new_n290_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1326gat));
  INV_X1    g465(.A(G22gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n636_), .B2(new_n511_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT42), .Z(new_n669_));
  NAND3_X1  g468(.A1(new_n645_), .A2(new_n667_), .A3(new_n511_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1327gat));
  NAND2_X1  g470(.A1(new_n579_), .A2(new_n583_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n635_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT108), .ZN(new_n674_));
  INV_X1    g473(.A(new_n622_), .ZN(new_n675_));
  NOR4_X1   g474(.A1(new_n516_), .A2(new_n674_), .A3(new_n640_), .A4(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n498_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n516_), .B2(new_n643_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n398_), .A2(new_n402_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n484_), .A2(new_n493_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n477_), .B1(new_n500_), .B2(new_n408_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .A4(new_n507_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n512_), .A2(new_n682_), .A3(new_n289_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n513_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n403_), .A3(new_n515_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n641_), .A2(new_n642_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n678_), .A2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n675_), .A2(new_n640_), .A3(new_n635_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(KEYINPUT105), .A3(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n687_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT43), .B(new_n643_), .C1(new_n683_), .C2(new_n685_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n691_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT44), .B(new_n691_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT107), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n690_), .A2(new_n702_), .A3(KEYINPUT44), .A4(new_n691_), .ZN(new_n703_));
  AOI22_X1  g502(.A1(new_n692_), .A2(new_n699_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n648_), .A2(G29gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n677_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n704_), .B2(new_n513_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n676_), .A2(new_n708_), .A3(new_n513_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT45), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n709_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n699_), .A2(new_n692_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n701_), .A2(new_n703_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n513_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G36gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(KEYINPUT46), .A3(new_n711_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n713_), .A2(new_n718_), .ZN(G1329gat));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(G43gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n704_), .B2(new_n290_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n676_), .A2(new_n721_), .A3(new_n290_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n714_), .A2(new_n290_), .A3(new_n715_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G43gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(KEYINPUT47), .A3(new_n723_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1330gat));
  AOI21_X1  g528(.A(G50gat), .B1(new_n676_), .B2(new_n511_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n511_), .A2(G50gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n704_), .B2(new_n731_), .ZN(G1331gat));
  AND4_X1   g531(.A1(new_n640_), .A2(new_n585_), .A3(new_n675_), .A4(new_n635_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n498_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n635_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n688_), .A2(new_n735_), .ZN(new_n736_));
  AND4_X1   g535(.A1(new_n686_), .A2(new_n736_), .A3(new_n640_), .A4(new_n675_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n648_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(G57gat), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n734_), .A2(G57gat), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT109), .Z(G1332gat));
  INV_X1    g540(.A(G64gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n733_), .B2(new_n513_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT48), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n737_), .A2(new_n742_), .A3(new_n513_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1333gat));
  AOI21_X1  g545(.A(new_n264_), .B1(new_n733_), .B2(new_n290_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT49), .Z(new_n748_));
  NOR2_X1   g547(.A1(new_n289_), .A2(G71gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT110), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n737_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n733_), .B2(new_n511_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT50), .Z(new_n755_));
  NAND2_X1  g554(.A1(new_n511_), .A2(new_n753_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT111), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n737_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1335gat));
  NOR4_X1   g558(.A1(new_n516_), .A2(new_n674_), .A3(new_n233_), .A4(new_n622_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n648_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n675_), .A2(new_n640_), .A3(new_n735_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT112), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n690_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n498_), .A2(G85gat), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT113), .Z(new_n766_));
  AOI21_X1  g565(.A(new_n761_), .B1(new_n764_), .B2(new_n766_), .ZN(G1336gat));
  AOI21_X1  g566(.A(G92gat), .B1(new_n760_), .B2(new_n513_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT114), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n513_), .A2(G92gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n764_), .B2(new_n770_), .ZN(G1337gat));
  AND3_X1   g570(.A1(new_n760_), .A2(new_n290_), .A3(new_n517_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n764_), .A2(new_n290_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(G99gat), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g574(.A1(new_n760_), .A2(new_n518_), .A3(new_n511_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n690_), .A2(new_n511_), .A3(new_n763_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(G106gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n736_), .A2(new_n783_), .A3(new_n640_), .A4(new_n622_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT54), .B1(new_n644_), .B2(new_n233_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n598_), .B(KEYINPUT12), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n596_), .A2(KEYINPUT66), .A3(new_n586_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(KEYINPUT55), .A3(new_n607_), .A4(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n586_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n601_), .A2(new_n603_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n596_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n789_), .A2(new_n792_), .A3(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n613_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n797_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n613_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n797_), .A2(new_n613_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n800_), .A2(new_n801_), .A3(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n213_), .B1(new_n221_), .B2(new_n209_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n217_), .B1(new_n806_), .B2(KEYINPUT116), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(KEYINPUT116), .B2(new_n806_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n229_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n230_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n616_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n787_), .B1(new_n805_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n800_), .A2(new_n801_), .A3(new_n804_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(KEYINPUT58), .A3(new_n616_), .A4(new_n813_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n815_), .B(new_n817_), .C1(new_n642_), .C2(new_n641_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n804_), .A2(new_n798_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n233_), .A2(new_n616_), .A3(KEYINPUT115), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT115), .B1(new_n233_), .B2(new_n616_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n822_), .A2(new_n825_), .B1(new_n617_), .B2(new_n813_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n821_), .B1(new_n826_), .B2(new_n584_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n798_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n797_), .B2(new_n613_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n813_), .A2(new_n617_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n672_), .A3(new_n820_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n827_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n818_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n735_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n786_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  NOR4_X1   g637(.A1(new_n738_), .A2(new_n511_), .A3(new_n513_), .A4(new_n289_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n818_), .A2(new_n834_), .A3(KEYINPUT120), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT120), .B1(new_n818_), .B2(new_n834_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n635_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n784_), .A2(new_n785_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT121), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n835_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n735_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n846_), .B(new_n786_), .C1(new_n849_), .C2(new_n841_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n845_), .A2(new_n850_), .A3(new_n839_), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n640_), .B(new_n840_), .C1(new_n851_), .C2(KEYINPUT59), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n233_), .A2(new_n272_), .ZN(new_n853_));
  OAI22_X1  g652(.A1(new_n852_), .A2(new_n272_), .B1(new_n851_), .B2(new_n853_), .ZN(G1340gat));
  INV_X1    g653(.A(new_n851_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n270_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n855_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n270_), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n622_), .B(new_n840_), .C1(new_n851_), .C2(KEYINPUT59), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n270_), .ZN(G1341gat));
  AOI211_X1 g658(.A(new_n735_), .B(new_n840_), .C1(new_n851_), .C2(KEYINPUT59), .ZN(new_n860_));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n635_), .A2(new_n861_), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n860_), .A2(new_n861_), .B1(new_n851_), .B2(new_n862_), .ZN(G1342gat));
  AOI21_X1  g662(.A(G134gat), .B1(new_n855_), .B2(new_n584_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n840_), .B1(new_n851_), .B2(KEYINPUT59), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT122), .B(G134gat), .Z(new_n866_));
  NOR2_X1   g665(.A1(new_n643_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n864_), .B1(new_n865_), .B2(new_n867_), .ZN(G1343gat));
  AND2_X1   g667(.A1(new_n845_), .A2(new_n850_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n684_), .A2(new_n511_), .A3(new_n289_), .A4(new_n648_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT123), .Z(new_n871_));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n233_), .A3(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n675_), .A3(new_n871_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g674(.A1(new_n869_), .A2(new_n635_), .A3(new_n871_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  NAND2_X1  g677(.A1(new_n869_), .A2(new_n871_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G162gat), .B1(new_n879_), .B2(new_n643_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n672_), .A2(G162gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n879_), .B2(new_n881_), .ZN(G1347gat));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n684_), .A2(new_n289_), .A3(new_n648_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n837_), .A2(new_n403_), .A3(new_n233_), .A4(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n416_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n885_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT62), .B1(new_n885_), .B2(G169gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n883_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n890_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n892_), .A2(new_n887_), .A3(KEYINPUT124), .A4(new_n888_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1348gat));
  AOI21_X1  g693(.A(new_n511_), .B1(new_n786_), .B2(new_n836_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n884_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n242_), .B1(new_n896_), .B2(new_n622_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n884_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n898_), .A2(new_n242_), .A3(new_n622_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n845_), .A2(new_n403_), .A3(new_n850_), .A4(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n897_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1349gat));
  NAND4_X1  g702(.A1(new_n869_), .A2(new_n403_), .A3(new_n635_), .A4(new_n884_), .ZN(new_n904_));
  INV_X1    g703(.A(G183gat), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n898_), .A2(new_n414_), .A3(new_n735_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n904_), .A2(new_n905_), .B1(new_n895_), .B2(new_n906_), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n896_), .B2(new_n643_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n584_), .A2(new_n251_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n896_), .B2(new_n909_), .ZN(G1351gat));
  NOR4_X1   g709(.A1(new_n684_), .A2(new_n403_), .A3(new_n498_), .A4(new_n290_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n845_), .A2(new_n233_), .A3(new_n850_), .A4(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(KEYINPUT126), .B2(new_n327_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT126), .B(G197gat), .Z(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n912_), .B2(new_n914_), .ZN(G1352gat));
  NAND3_X1  g714(.A1(new_n869_), .A2(new_n675_), .A3(new_n911_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g716(.A1(new_n845_), .A2(new_n635_), .A3(new_n850_), .A4(new_n911_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  AND2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n918_), .B2(new_n919_), .ZN(G1354gat));
  NAND4_X1  g721(.A1(new_n845_), .A2(new_n688_), .A3(new_n850_), .A4(new_n911_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(G218gat), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n672_), .A2(G218gat), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n845_), .A2(new_n850_), .A3(new_n911_), .A4(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n924_), .A2(KEYINPUT127), .A3(new_n926_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1355gat));
endmodule


