//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G197gat), .A2(G204gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT85), .B(G204gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n203_), .B1(new_n204_), .B2(G197gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  NOR3_X1   g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT87), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT86), .ZN(new_n211_));
  INV_X1    g010(.A(G197gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n211_), .B(new_n212_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT21), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT86), .B1(new_n212_), .B2(G204gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(new_n204_), .B2(new_n212_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n210_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n217_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n222_), .A2(KEYINPUT87), .A3(KEYINPUT21), .A4(new_n215_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n208_), .B1(new_n205_), .B2(KEYINPUT21), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n209_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G183gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT25), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G183gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT78), .B(G190gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT26), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n229_), .B(new_n231_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G169gat), .ZN(new_n237_));
  INV_X1    g036(.A(G176gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n240_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n242_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n232_), .A2(new_n228_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n247_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT22), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n238_), .B1(new_n255_), .B2(KEYINPUT79), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(new_n237_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n236_), .A2(new_n249_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT93), .B1(new_n227_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT93), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n225_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n260_), .B(new_n261_), .C1(new_n262_), .C2(new_n209_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT20), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT90), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n229_), .A2(new_n231_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n268_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G190gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n242_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n248_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n237_), .A2(KEYINPUT22), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n255_), .A2(G169gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n238_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n239_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(KEYINPUT92), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT92), .ZN(new_n283_));
  OR2_X1    g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n282_), .A2(new_n283_), .B1(new_n253_), .B2(new_n284_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n274_), .A2(new_n276_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n286_));
  AOI211_X1 g085(.A(new_n265_), .B(new_n267_), .C1(new_n227_), .C2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n224_), .A2(new_n226_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n209_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n258_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n242_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n229_), .A2(new_n231_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT90), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n273_), .A3(new_n269_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT91), .B1(new_n253_), .B2(new_n243_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n248_), .A2(new_n275_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n291_), .B(new_n294_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n285_), .A2(new_n281_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n262_), .B2(new_n209_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n290_), .A2(new_n300_), .A3(KEYINPUT20), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n264_), .A2(new_n287_), .B1(new_n301_), .B2(new_n267_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G8gat), .B(G36gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n202_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n264_), .A2(new_n287_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n301_), .A2(new_n267_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n307_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n202_), .A3(new_n312_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(G228gat), .A2(G233gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n227_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(KEYINPUT1), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(G155gat), .B2(G162gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n327_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n328_), .B1(new_n331_), .B2(KEYINPUT81), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n333_), .A3(new_n327_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n326_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n324_), .A2(KEYINPUT82), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n322_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340_));
  OAI22_X1  g139(.A1(new_n340_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n337_), .A2(new_n339_), .A3(new_n341_), .A4(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n327_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n321_), .B1(new_n335_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G155gat), .ZN(new_n350_));
  INV_X1    g149(.A(G162gat), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT1), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT81), .B1(new_n352_), .B2(new_n344_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n328_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n334_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n325_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(KEYINPUT83), .A3(new_n347_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n349_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n319_), .B1(new_n320_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT88), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n355_), .A2(new_n325_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(new_n320_), .ZN(new_n362_));
  OAI211_X1 g161(.A(KEYINPUT88), .B(KEYINPUT29), .C1(new_n335_), .C2(new_n348_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n362_), .B(new_n363_), .C1(new_n262_), .C2(new_n209_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n364_), .A2(KEYINPUT89), .A3(new_n318_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT89), .B1(new_n364_), .B2(new_n318_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n359_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G78gat), .B(G106gat), .Z(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G22gat), .B(G50gat), .Z(new_n370_));
  XOR2_X1   g169(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n358_), .A2(new_n320_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n372_), .B1(new_n358_), .B2(new_n320_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n370_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n370_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n373_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n368_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n382_), .B(new_n359_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n369_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n364_), .A2(new_n318_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n364_), .A2(KEYINPUT89), .A3(new_n318_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n382_), .B1(new_n389_), .B2(new_n359_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n383_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n380_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n315_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n267_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n265_), .B1(new_n227_), .B2(new_n286_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n264_), .B2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n301_), .A2(new_n267_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n393_), .B1(new_n307_), .B2(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n317_), .A2(new_n384_), .A3(new_n392_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT100), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n369_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n381_), .B1(new_n369_), .B2(new_n383_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT100), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n317_), .A4(new_n399_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT80), .B(G15gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n258_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G127gat), .B(G134gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G113gat), .B(G120gat), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n413_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n411_), .B(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G71gat), .B(G99gat), .Z(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(G43gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT30), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT31), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n418_), .B(new_n422_), .Z(new_n423_));
  NAND3_X1  g222(.A1(new_n349_), .A2(new_n357_), .A3(new_n417_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(KEYINPUT96), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n416_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n361_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n428_), .A3(KEYINPUT4), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT97), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n424_), .A2(new_n428_), .A3(KEYINPUT97), .A4(KEYINPUT4), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n349_), .A2(new_n357_), .A3(new_n434_), .A4(new_n417_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n436_), .B(KEYINPUT98), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n424_), .A2(new_n428_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(new_n437_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G29gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G85gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT0), .B(G57gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  NAND3_X1  g246(.A1(new_n440_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n438_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n449_), .B1(new_n450_), .B2(new_n442_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n423_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n392_), .A2(new_n384_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n452_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n317_), .A4(new_n399_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n437_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n449_), .B1(new_n441_), .B2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n435_), .A2(new_n457_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n433_), .B2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n442_), .B1(new_n433_), .B2(new_n439_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT33), .B1(new_n462_), .B2(new_n447_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464_));
  NOR4_X1   g263(.A1(new_n450_), .A2(new_n464_), .A3(new_n442_), .A4(new_n449_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT99), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n307_), .A2(KEYINPUT32), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n398_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  OAI211_X1 g269(.A(KEYINPUT99), .B(new_n470_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n448_), .A2(new_n451_), .B1(new_n468_), .B2(new_n302_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n461_), .A2(new_n466_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n456_), .B1(new_n474_), .B2(new_n454_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n407_), .A2(new_n453_), .B1(new_n475_), .B2(new_n423_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G230gat), .A2(G233gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT6), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n480_));
  OR3_X1    g279(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G85gat), .B(G92gat), .Z(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT65), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT8), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n482_), .B(new_n483_), .C1(new_n485_), .C2(KEYINPUT8), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(KEYINPUT9), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT10), .B(G99gat), .Z(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT64), .B(G92gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT9), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(G85gat), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n489_), .A2(new_n492_), .A3(new_n479_), .A4(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n487_), .A2(new_n488_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n499_));
  XOR2_X1   g298(.A(G71gat), .B(G78gat), .Z(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n499_), .A2(new_n500_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n497_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(new_n504_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n477_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT66), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT67), .B1(new_n497_), .B2(new_n504_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT12), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n511_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n512_), .A2(new_n477_), .A3(new_n513_), .A4(new_n505_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(new_n508_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G120gat), .B(G148gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT5), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G176gat), .B(G204gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n509_), .A2(new_n514_), .A3(new_n515_), .A4(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n507_), .B(KEYINPUT66), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n524_), .A2(KEYINPUT68), .A3(new_n514_), .A4(new_n520_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n514_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n519_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n526_), .A2(KEYINPUT13), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT13), .B1(new_n526_), .B2(new_n528_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G29gat), .B(G36gat), .Z(new_n532_));
  XOR2_X1   g331(.A(G43gat), .B(G50gat), .Z(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT15), .Z(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT74), .B(G8gat), .Z(new_n536_));
  INV_X1    g335(.A(G1gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT14), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G8gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n535_), .A2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n534_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n545_), .B(new_n534_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n550_), .B1(new_n551_), .B2(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT77), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G169gat), .B(G197gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n553_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n531_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n476_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n560_), .A2(KEYINPUT37), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(KEYINPUT37), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n535_), .A2(new_n497_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT35), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(KEYINPUT35), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT70), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n569_), .B2(KEYINPUT72), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n563_), .B(new_n570_), .C1(new_n497_), .C2(new_n534_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(KEYINPUT72), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n572_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT71), .ZN(new_n576_));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT36), .Z(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n574_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n578_), .A2(KEYINPUT36), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n561_), .B(new_n562_), .C1(new_n581_), .C2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n586_), .A2(new_n560_), .A3(KEYINPUT37), .A4(new_n580_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n504_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(new_n545_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G127gat), .B(G155gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT17), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n596_), .A2(KEYINPUT17), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n591_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n588_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT76), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n559_), .A2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n605_), .A2(G1gat), .A3(new_n455_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(KEYINPUT38), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(KEYINPUT38), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n581_), .A2(new_n584_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n476_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n558_), .A2(new_n602_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G1gat), .B1(new_n612_), .B2(new_n455_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n607_), .A2(new_n608_), .A3(new_n613_), .ZN(G1324gat));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n317_), .A2(new_n399_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G8gat), .B1(new_n612_), .B2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n615_), .B1(new_n618_), .B2(KEYINPUT101), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(KEYINPUT101), .B2(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(KEYINPUT101), .A3(new_n615_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n559_), .A2(new_n536_), .A3(new_n604_), .A4(new_n616_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n620_), .A2(KEYINPUT40), .A3(new_n621_), .A4(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1325gat));
  OAI21_X1  g426(.A(G15gat), .B1(new_n612_), .B2(new_n423_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT41), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n605_), .A2(G15gat), .A3(new_n423_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1326gat));
  OAI21_X1  g430(.A(G22gat), .B1(new_n612_), .B2(new_n404_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT42), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n404_), .A2(G22gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n633_), .B1(new_n605_), .B2(new_n634_), .ZN(G1327gat));
  NAND2_X1  g434(.A1(new_n407_), .A2(new_n453_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n461_), .A2(new_n466_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n472_), .A2(new_n473_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n454_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n455_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n616_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n423_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n636_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n609_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n601_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n643_), .A2(new_n531_), .A3(new_n557_), .A4(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G29gat), .B1(new_n647_), .B2(new_n452_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n558_), .A2(new_n601_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n588_), .B(KEYINPUT102), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT43), .B1(new_n476_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n643_), .A2(new_n654_), .A3(new_n588_), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n649_), .B(new_n651_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n588_), .B(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n643_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n588_), .A2(new_n654_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n476_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n650_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT44), .B1(new_n662_), .B2(KEYINPUT103), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n651_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n656_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n452_), .A2(G29gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n648_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n667_), .B2(new_n616_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n616_), .A2(new_n671_), .ZN(new_n673_));
  OR3_X1    g472(.A1(new_n646_), .A2(KEYINPUT104), .A3(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT104), .B1(new_n646_), .B2(new_n673_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(KEYINPUT45), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n670_), .B1(new_n672_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n664_), .A2(KEYINPUT44), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n649_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT103), .B(new_n651_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G36gat), .B1(new_n685_), .B2(new_n617_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n678_), .A2(new_n679_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(KEYINPUT46), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n681_), .A2(new_n688_), .ZN(G1329gat));
  XOR2_X1   g488(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n423_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n692_), .B(new_n682_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G43gat), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n646_), .A2(G43gat), .A3(new_n423_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n691_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n690_), .B(new_n695_), .C1(new_n693_), .C2(G43gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1330gat));
  INV_X1    g498(.A(G50gat), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n404_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n667_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n646_), .B2(new_n404_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n702_), .A2(KEYINPUT106), .A3(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1331gat));
  INV_X1    g507(.A(new_n557_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n601_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n531_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n610_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(G57gat), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n455_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n476_), .A2(new_n531_), .A3(new_n557_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n604_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n455_), .B1(new_n716_), .B2(KEYINPUT107), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(KEYINPUT107), .B2(new_n716_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n718_), .B2(new_n713_), .ZN(G1332gat));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720_));
  INV_X1    g519(.A(new_n712_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n616_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(G64gat), .ZN(new_n723_));
  INV_X1    g522(.A(G64gat), .ZN(new_n724_));
  AOI211_X1 g523(.A(KEYINPUT48), .B(new_n724_), .C1(new_n721_), .C2(new_n616_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n616_), .A2(new_n724_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT108), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n723_), .A2(new_n725_), .B1(new_n716_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT109), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n712_), .B2(new_n423_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT49), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n423_), .A2(G71gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n716_), .B2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n712_), .B2(new_n404_), .ZN(new_n734_));
  XOR2_X1   g533(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n404_), .A2(G78gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n716_), .B2(new_n737_), .ZN(G1335gat));
  AND2_X1   g537(.A1(new_n715_), .A2(new_n645_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n452_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n653_), .A2(new_n655_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n531_), .A2(new_n601_), .A3(new_n557_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT111), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n452_), .A2(G85gat), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT112), .Z(new_n746_));
  AOI21_X1  g545(.A(new_n740_), .B1(new_n744_), .B2(new_n746_), .ZN(G1336gat));
  AOI21_X1  g546(.A(G92gat), .B1(new_n739_), .B2(new_n616_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n616_), .A2(new_n493_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n744_), .B2(new_n749_), .ZN(G1337gat));
  NAND2_X1  g549(.A1(new_n744_), .A2(new_n692_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n692_), .A2(new_n490_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n751_), .A2(G99gat), .B1(new_n739_), .B2(new_n752_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g553(.A1(new_n739_), .A2(new_n491_), .A3(new_n454_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n741_), .A2(new_n454_), .A3(new_n743_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G106gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G106gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g560(.A(new_n513_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n505_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n763_));
  OAI211_X1 g562(.A(G230gat), .B(G233gat), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n514_), .A3(KEYINPUT55), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n762_), .A2(new_n763_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n477_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n765_), .A2(KEYINPUT113), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT113), .B1(new_n765_), .B2(new_n768_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n519_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n557_), .A2(new_n526_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n519_), .B(new_n772_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n526_), .A2(new_n528_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n552_), .A2(new_n556_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n549_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n547_), .A2(new_n548_), .A3(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n551_), .A2(new_n781_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n556_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n779_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n609_), .B1(new_n778_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n771_), .A2(KEYINPUT56), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(KEYINPUT58), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n519_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n526_), .A2(new_n785_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n788_), .A2(new_n791_), .A3(new_n793_), .A4(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n588_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n765_), .A2(new_n768_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n765_), .A2(KEYINPUT113), .A3(new_n768_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n520_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n794_), .B1(new_n802_), .B2(new_n792_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n791_), .B1(new_n803_), .B2(new_n788_), .ZN(new_n804_));
  OAI22_X1  g603(.A1(new_n787_), .A2(KEYINPUT57), .B1(new_n797_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n775_), .B1(new_n802_), .B2(new_n772_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n806_), .A2(new_n774_), .B1(new_n779_), .B2(new_n785_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n609_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n602_), .B1(new_n805_), .B2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n588_), .A2(new_n710_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n531_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(new_n531_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n810_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n407_), .A2(new_n452_), .A3(new_n692_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT116), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G113gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n557_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(KEYINPUT59), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n709_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n827_), .B2(new_n822_), .ZN(G1340gat));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n531_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n821_), .B(new_n830_), .C1(KEYINPUT60), .C2(new_n829_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n531_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n829_), .ZN(G1341gat));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n821_), .A2(new_n834_), .A3(new_n601_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n602_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n834_), .ZN(G1342gat));
  NAND2_X1  g636(.A1(new_n824_), .A2(new_n826_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n588_), .ZN(new_n839_));
  INV_X1    g638(.A(G134gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n820_), .B2(new_n644_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT117), .B(new_n840_), .C1(new_n820_), .C2(new_n644_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n838_), .A2(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(G1343gat));
  NAND3_X1  g645(.A1(new_n454_), .A2(new_n452_), .A3(new_n423_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n616_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n817_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n709_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT118), .B(G141gat), .Z(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1344gat));
  OAI21_X1  g651(.A(new_n808_), .B1(new_n807_), .B2(new_n609_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n787_), .A2(KEYINPUT57), .ZN(new_n854_));
  INV_X1    g653(.A(new_n788_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n795_), .A2(new_n793_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n790_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(new_n588_), .A3(new_n796_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n853_), .A2(new_n854_), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n815_), .B1(new_n859_), .B2(new_n602_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n860_), .A2(new_n616_), .A3(new_n847_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n529_), .A2(new_n530_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n861_), .A2(new_n865_), .A3(new_n601_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT119), .B1(new_n849_), .B2(new_n602_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1346gat));
  AOI21_X1  g670(.A(G162gat), .B1(new_n861_), .B2(new_n609_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n849_), .A2(new_n351_), .A3(new_n652_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1347gat));
  NAND3_X1  g673(.A1(new_n616_), .A2(new_n404_), .A3(new_n453_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n810_), .B2(new_n816_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n557_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT121), .Z(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  INV_X1    g679(.A(new_n875_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n817_), .A2(KEYINPUT120), .A3(new_n557_), .A4(new_n881_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(G169gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT120), .B1(new_n876_), .B2(new_n557_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n880_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(G169gat), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n887_), .A2(KEYINPUT62), .A3(new_n884_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n879_), .B1(new_n886_), .B2(new_n888_), .ZN(G1348gat));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  INV_X1    g689(.A(new_n876_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n531_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n892_), .B2(G176gat), .ZN(new_n893_));
  OAI211_X1 g692(.A(KEYINPUT122), .B(new_n238_), .C1(new_n891_), .C2(new_n531_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n876_), .A2(G176gat), .A3(new_n862_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n896_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n893_), .A2(new_n894_), .B1(new_n897_), .B2(new_n898_), .ZN(G1349gat));
  NAND2_X1  g698(.A1(new_n876_), .A2(new_n601_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n272_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n228_), .B2(new_n900_), .ZN(G1350gat));
  OAI21_X1  g701(.A(G190gat), .B1(new_n891_), .B2(new_n839_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n876_), .A2(new_n609_), .A3(new_n273_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1351gat));
  NAND3_X1  g704(.A1(new_n454_), .A2(new_n455_), .A3(new_n423_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n907_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n908_), .A2(new_n616_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n860_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n557_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g713(.A(G204gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n817_), .A2(new_n910_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n531_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n912_), .A2(new_n204_), .A3(new_n862_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1353gat));
  NAND2_X1  g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n601_), .A2(new_n922_), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT126), .Z(new_n924_));
  NOR3_X1   g723(.A1(new_n916_), .A2(KEYINPUT127), .A3(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926_));
  INV_X1    g725(.A(new_n924_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n912_), .B2(new_n927_), .ZN(new_n928_));
  OR2_X1    g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  OR3_X1    g728(.A1(new_n925_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n925_), .B2(new_n928_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1354gat));
  OR3_X1    g731(.A1(new_n916_), .A2(G218gat), .A3(new_n644_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G218gat), .B1(new_n916_), .B2(new_n839_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1355gat));
endmodule


