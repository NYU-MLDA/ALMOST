//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(G92gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n203_), .A2(new_n206_), .A3(new_n208_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT7), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n214_), .A2(new_n218_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT68), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n214_), .A2(new_n218_), .ZN(new_n223_));
  AND2_X1   g022(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n222_), .B(new_n223_), .C1(new_n226_), .C2(new_n214_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n221_), .A2(new_n208_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n202_), .A2(KEYINPUT67), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G85gat), .B(G92gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n213_), .B1(new_n228_), .B2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n213_), .A3(new_n232_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n219_), .A2(new_n220_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n208_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n212_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G29gat), .B(G36gat), .Z(new_n239_));
  XOR2_X1   g038(.A(G43gat), .B(G50gat), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT15), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n238_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G232gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n245_), .ZN(new_n251_));
  OAI221_X1 g050(.A(new_n247_), .B1(KEYINPUT35), .B2(new_n250_), .C1(new_n238_), .C2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(KEYINPUT35), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G190gat), .B(G218gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G134gat), .B(G162gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT36), .Z(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n257_), .A2(KEYINPUT36), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT37), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT37), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n260_), .A2(new_n265_), .A3(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G57gat), .B(G64gat), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT11), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(KEYINPUT11), .ZN(new_n270_));
  XOR2_X1   g069(.A(G71gat), .B(G78gat), .Z(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n270_), .A2(new_n271_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G231gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT71), .B(G8gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G1gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT14), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G15gat), .B(G22gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G8gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n276_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G127gat), .B(G155gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G183gat), .B(G211gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT17), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n286_), .A2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n291_), .A2(KEYINPUT17), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n286_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n267_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT73), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n300_));
  INV_X1    g099(.A(new_n274_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n238_), .A2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n274_), .B(new_n212_), .C1(new_n234_), .C2(new_n237_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT12), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT12), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n238_), .A2(new_n305_), .A3(new_n301_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G230gat), .A2(G233gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT64), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n302_), .A2(new_n303_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n309_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G120gat), .B(G148gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT5), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G176gat), .B(G204gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n318_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n311_), .A2(new_n313_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT13), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n319_), .A2(KEYINPUT13), .A3(new_n321_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT69), .Z(new_n327_));
  OR3_X1    g126(.A1(new_n299_), .A2(new_n300_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329_));
  XOR2_X1   g128(.A(G8gat), .B(G36gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT81), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT80), .B1(new_n341_), .B2(G190gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT25), .B(G183gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(G190gat), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n342_), .B(new_n343_), .C1(new_n344_), .C2(KEYINPUT80), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n337_), .B(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n340_), .B(new_n345_), .C1(new_n349_), .C2(new_n339_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G183gat), .A3(G190gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT82), .ZN(new_n353_));
  INV_X1    g152(.A(G183gat), .ZN(new_n354_));
  INV_X1    g153(.A(G190gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT23), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n350_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(KEYINPUT83), .B(G176gat), .Z(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT22), .B(G169gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n356_), .A2(new_n352_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n361_), .B(new_n348_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G197gat), .B(G204gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT21), .ZN(new_n368_));
  OR3_X1    g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n366_), .A2(new_n368_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n368_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n367_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n369_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n336_), .B1(new_n365_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n348_), .B(KEYINPUT92), .Z(new_n379_));
  OAI211_X1 g178(.A(new_n361_), .B(new_n379_), .C1(new_n357_), .C2(new_n363_), .ZN(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n381_));
  AOI21_X1  g180(.A(new_n362_), .B1(new_n337_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n344_), .A2(new_n343_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n382_), .B(new_n383_), .C1(new_n349_), .C2(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n385_), .A2(new_n373_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n374_), .A2(new_n378_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT20), .B1(new_n365_), .B2(new_n373_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT90), .B(KEYINPUT20), .C1(new_n365_), .C2(new_n373_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n385_), .A2(KEYINPUT93), .A3(new_n373_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n385_), .A2(new_n373_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT93), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .A4(new_n396_), .ZN(new_n397_));
  AOI211_X1 g196(.A(new_n335_), .B(new_n388_), .C1(new_n397_), .C2(new_n377_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n391_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n392_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n377_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n334_), .B1(new_n401_), .B2(new_n387_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n329_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G71gat), .B(G99gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT84), .B(G43gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(G15gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT30), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n358_), .B2(new_n364_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n358_), .A2(new_n364_), .A3(new_n410_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n407_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n415_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G127gat), .B(G134gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT85), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n419_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT31), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT86), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(KEYINPUT86), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G22gat), .B(G50gat), .ZN(new_n429_));
  INV_X1    g228(.A(G228gat), .ZN(new_n430_));
  INV_X1    g229(.A(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT88), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n373_), .B(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n434_), .A2(KEYINPUT1), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G155gat), .A2(G162gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n436_), .B2(KEYINPUT1), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT87), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n435_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n438_), .B2(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G141gat), .A2(G148gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n440_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n436_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n434_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n442_), .B(KEYINPUT3), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n441_), .B(KEYINPUT2), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT29), .B1(new_n444_), .B2(new_n449_), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n430_), .B(new_n431_), .C1(new_n433_), .C2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n373_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n429_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n454_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n433_), .A2(new_n450_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(G228gat), .A3(G233gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n429_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT28), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n444_), .A2(new_n449_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G78gat), .B(G106gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n466_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n467_), .B1(new_n470_), .B2(new_n464_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n455_), .A2(new_n460_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n455_), .A2(new_n460_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n428_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n455_), .A2(new_n460_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n469_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n478_), .A2(new_n425_), .A3(new_n427_), .A4(new_n472_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT4), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n444_), .A2(new_n449_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n422_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT95), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n419_), .B(new_n420_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n462_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n486_), .A3(new_n422_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n483_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n462_), .A2(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n483_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n482_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G1gat), .B(G29gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G57gat), .B(G85gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  NAND3_X1  g299(.A1(new_n489_), .A2(new_n481_), .A3(new_n490_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n495_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n500_), .B1(new_n495_), .B2(new_n501_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n374_), .B1(new_n385_), .B2(new_n433_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n377_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n397_), .B2(new_n377_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n335_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n388_), .B1(new_n397_), .B2(new_n377_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n334_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n511_), .A3(KEYINPUT27), .ZN(new_n512_));
  AND4_X1   g311(.A1(new_n403_), .A2(new_n480_), .A3(new_n505_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n504_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n502_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n508_), .A2(KEYINPUT32), .A3(new_n334_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n510_), .B1(new_n517_), .B2(new_n335_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT97), .B1(new_n504_), .B2(KEYINPUT33), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n398_), .A2(new_n402_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n504_), .A2(KEYINPUT33), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n491_), .A2(new_n482_), .A3(new_n494_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n489_), .A2(new_n490_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n482_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n500_), .A3(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .A4(new_n526_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n504_), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n519_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n478_), .A2(new_n472_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(new_n428_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n513_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT75), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n245_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n285_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n251_), .A2(KEYINPUT75), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n245_), .A2(new_n536_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n539_), .B(new_n540_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n541_), .A3(KEYINPUT76), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT76), .B1(new_n538_), .B2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n535_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n285_), .A2(new_n246_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n546_), .A2(new_n541_), .A3(new_n547_), .A4(new_n534_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n541_), .A3(new_n534_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT77), .ZN(new_n550_));
  XOR2_X1   g349(.A(G113gat), .B(G141gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT78), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G169gat), .B(G197gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n552_), .B(new_n553_), .Z(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n545_), .A2(new_n548_), .A3(new_n550_), .A4(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n538_), .A2(new_n541_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n534_), .B1(new_n559_), .B2(new_n542_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n550_), .A2(new_n548_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n554_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT79), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n556_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(KEYINPUT79), .B(new_n554_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n533_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n328_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n300_), .B1(new_n299_), .B2(new_n327_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n515_), .B(KEYINPUT98), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(G1gat), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(KEYINPUT38), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n529_), .A2(new_n532_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n513_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n326_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n578_), .A2(new_n296_), .A3(new_n566_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n263_), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G1gat), .B1(new_n580_), .B2(new_n505_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582_));
  INV_X1    g381(.A(new_n573_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n582_), .B1(new_n570_), .B2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n574_), .A2(new_n581_), .A3(new_n584_), .ZN(G1324gat));
  NAND2_X1  g384(.A1(new_n403_), .A2(new_n512_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(G8gat), .B1(new_n580_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT99), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(KEYINPUT39), .A3(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(KEYINPUT39), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n587_), .A2(new_n277_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n328_), .A2(new_n569_), .A3(new_n567_), .A4(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT40), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n592_), .A2(new_n593_), .A3(KEYINPUT40), .A4(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(G1325gat));
  INV_X1    g399(.A(new_n428_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(G15gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n571_), .A2(KEYINPUT100), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G15gat), .B1(new_n580_), .B2(new_n601_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT41), .Z(new_n605_));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606_));
  INV_X1    g405(.A(new_n602_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n606_), .B1(new_n570_), .B2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n603_), .A2(new_n605_), .A3(new_n608_), .ZN(G1326gat));
  OAI21_X1  g408(.A(G22gat), .B1(new_n580_), .B2(new_n530_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT42), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n530_), .A2(G22gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n611_), .B1(new_n570_), .B2(new_n612_), .ZN(G1327gat));
  INV_X1    g412(.A(new_n263_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n296_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT102), .B1(new_n263_), .B2(new_n297_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n578_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n567_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(G29gat), .B1(new_n620_), .B2(new_n515_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT43), .B1(new_n533_), .B2(new_n267_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT43), .ZN(new_n623_));
  INV_X1    g422(.A(new_n267_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n532_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n528_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n402_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n627_), .A2(new_n526_), .A3(new_n511_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n626_), .A2(new_n628_), .A3(new_n520_), .A4(new_n522_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n625_), .B1(new_n629_), .B2(new_n519_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n623_), .B(new_n624_), .C1(new_n630_), .C2(new_n513_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n622_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n564_), .A2(new_n565_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n326_), .A2(new_n296_), .A3(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT101), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(KEYINPUT44), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT44), .B1(new_n632_), .B2(new_n635_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n572_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(G29gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n621_), .B1(new_n639_), .B2(new_n641_), .ZN(G1328gat));
  NOR2_X1   g441(.A1(new_n587_), .A2(G36gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT45), .B1(new_n619_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT45), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n567_), .A2(new_n646_), .A3(new_n618_), .A4(new_n643_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n632_), .A2(new_n635_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n586_), .A3(new_n636_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n648_), .B1(new_n652_), .B2(G36gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n654_), .ZN(new_n656_));
  AOI211_X1 g455(.A(new_n656_), .B(new_n648_), .C1(new_n652_), .C2(G36gat), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1329gat));
  INV_X1    g457(.A(G43gat), .ZN(new_n659_));
  NOR4_X1   g458(.A1(new_n637_), .A2(new_n638_), .A3(new_n659_), .A4(new_n601_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n619_), .B2(new_n601_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(new_n662_), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT47), .B1(new_n660_), .B2(new_n665_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1330gat));
  AOI21_X1  g468(.A(G50gat), .B1(new_n620_), .B2(new_n531_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n531_), .A2(G50gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n639_), .B2(new_n671_), .ZN(G1331gat));
  NAND2_X1  g471(.A1(new_n577_), .A2(new_n263_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n327_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n566_), .A2(new_n297_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G57gat), .B1(new_n677_), .B2(new_n505_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n577_), .A2(new_n566_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n679_), .A2(new_n299_), .A3(new_n326_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n572_), .A2(G57gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1332gat));
  OAI21_X1  g481(.A(G64gat), .B1(new_n677_), .B2(new_n587_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT48), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n587_), .A2(G64gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n680_), .B2(new_n685_), .ZN(G1333gat));
  OR3_X1    g485(.A1(new_n680_), .A2(G71gat), .A3(new_n601_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n676_), .A2(new_n428_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT105), .B(KEYINPUT49), .Z(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(G71gat), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(G71gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1334gat));
  OAI21_X1  g491(.A(G78gat), .B1(new_n677_), .B2(new_n530_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n530_), .A2(G78gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n680_), .B2(new_n696_), .ZN(G1335gat));
  AND2_X1   g496(.A1(new_n616_), .A2(new_n617_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n679_), .A2(new_n674_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G85gat), .B1(new_n699_), .B2(new_n640_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n578_), .A2(new_n296_), .A3(new_n566_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n622_), .B2(new_n631_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(KEYINPUT107), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n705_), .B(new_n701_), .C1(new_n622_), .C2(new_n631_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n515_), .A2(new_n209_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n700_), .B1(new_n708_), .B2(new_n709_), .ZN(G1336gat));
  INV_X1    g509(.A(G92gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n699_), .A2(new_n711_), .A3(new_n586_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n587_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n711_), .ZN(G1337gat));
  AND3_X1   g513(.A1(new_n699_), .A2(new_n204_), .A3(new_n428_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n428_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(G99gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n718_), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n720_), .B(new_n715_), .C1(new_n716_), .C2(G99gat), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1338gat));
  AOI211_X1 g521(.A(new_n530_), .B(new_n701_), .C1(new_n622_), .C2(new_n631_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT109), .B1(new_n723_), .B2(new_n205_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n702_), .A2(new_n531_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(G106gat), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n724_), .A2(new_n727_), .A3(KEYINPUT52), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT109), .B(new_n729_), .C1(new_n723_), .C2(new_n205_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n699_), .A2(new_n205_), .A3(new_n531_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT53), .B1(new_n728_), .B2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n727_), .A3(KEYINPUT52), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n734_), .A2(new_n730_), .A3(new_n735_), .A4(new_n731_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(G1339gat));
  AOI21_X1  g536(.A(KEYINPUT110), .B1(new_n566_), .B2(new_n297_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n566_), .A2(new_n297_), .A3(KEYINPUT110), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n326_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n267_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n740_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(new_n738_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT111), .B1(new_n745_), .B2(new_n326_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT54), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n741_), .A2(new_n742_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(KEYINPUT111), .A3(new_n326_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT54), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .A4(new_n267_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n747_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n304_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n304_), .A2(KEYINPUT112), .A3(new_n309_), .A4(new_n306_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT55), .B1(new_n307_), .B2(new_n310_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759_));
  AOI211_X1 g558(.A(new_n759_), .B(new_n309_), .C1(new_n304_), .C2(new_n306_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n757_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT56), .B1(new_n761_), .B2(new_n320_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n311_), .A2(new_n759_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n307_), .A2(KEYINPUT55), .A3(new_n310_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n755_), .A4(new_n756_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n318_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n762_), .A2(new_n321_), .A3(new_n633_), .A4(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n321_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n765_), .A2(new_n318_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(KEYINPUT56), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n773_), .A2(KEYINPUT113), .A3(new_n633_), .A4(new_n767_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n534_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n546_), .A2(new_n541_), .A3(new_n535_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n554_), .A3(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n556_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n322_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n770_), .A2(new_n774_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n614_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n779_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n614_), .B1(new_n785_), .B2(new_n774_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n762_), .A2(new_n321_), .A3(new_n778_), .A4(new_n767_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT58), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n773_), .A2(new_n789_), .A3(new_n778_), .A4(new_n767_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT114), .B1(new_n791_), .B2(new_n624_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n793_), .B(new_n267_), .C1(new_n788_), .C2(new_n790_), .ZN(new_n794_));
  OAI221_X1 g593(.A(new_n783_), .B1(new_n786_), .B2(KEYINPUT57), .C1(new_n792_), .C2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n752_), .B1(new_n795_), .B2(new_n296_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n586_), .A2(new_n475_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n572_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT59), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n747_), .A2(new_n751_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n780_), .A2(new_n263_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n781_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n780_), .A2(new_n782_), .B1(new_n791_), .B2(new_n624_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n297_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n806_), .B2(KEYINPUT115), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n808_), .B(new_n297_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n801_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n800_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811_), .B2(new_n566_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n791_), .A2(new_n624_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n793_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n791_), .A2(KEYINPUT114), .A3(new_n624_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n803_), .A2(new_n781_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n297_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n798_), .B1(new_n818_), .B2(new_n752_), .ZN(new_n819_));
  OR3_X1    g618(.A1(new_n819_), .A2(G113gat), .A3(new_n566_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n812_), .A2(new_n820_), .ZN(G1340gat));
  XNOR2_X1  g620(.A(KEYINPUT116), .B(G120gat), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT60), .B1(new_n578_), .B2(new_n822_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n327_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n811_), .B2(new_n825_), .ZN(new_n826_));
  OR3_X1    g625(.A1(new_n819_), .A2(KEYINPUT60), .A3(new_n824_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(G1341gat));
  OAI21_X1  g627(.A(G127gat), .B1(new_n811_), .B2(new_n296_), .ZN(new_n829_));
  OR3_X1    g628(.A1(new_n819_), .A2(G127gat), .A3(new_n296_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1342gat));
  INV_X1    g630(.A(G134gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n819_), .B2(new_n263_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT117), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n835_), .B(new_n832_), .C1(new_n819_), .C2(new_n263_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n783_), .A2(new_n813_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n786_), .A2(KEYINPUT57), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n296_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n752_), .B1(new_n839_), .B2(new_n808_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n806_), .A2(KEYINPUT115), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n842_), .A2(new_n801_), .B1(new_n819_), .B2(KEYINPUT59), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n267_), .A2(new_n832_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n834_), .A2(new_n836_), .B1(new_n843_), .B2(new_n844_), .ZN(G1343gat));
  NOR2_X1   g644(.A1(new_n792_), .A2(new_n794_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n783_), .B1(new_n786_), .B2(KEYINPUT57), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n296_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n802_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n572_), .A2(new_n586_), .A3(new_n479_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(KEYINPUT118), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n566_), .ZN(new_n853_));
  XOR2_X1   g652(.A(KEYINPUT119), .B(G141gat), .Z(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1344gat));
  NOR2_X1   g654(.A1(new_n852_), .A2(new_n674_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT120), .B(G148gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1345gat));
  OAI211_X1 g657(.A(new_n297_), .B(new_n851_), .C1(new_n818_), .C2(new_n752_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT121), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n849_), .A2(new_n861_), .A3(new_n297_), .A4(new_n851_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n860_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1346gat));
  OAI21_X1  g665(.A(G162gat), .B1(new_n852_), .B2(new_n267_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n263_), .A2(G162gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n852_), .B2(new_n868_), .ZN(G1347gat));
  NAND2_X1  g668(.A1(new_n572_), .A2(new_n586_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n870_), .A2(new_n601_), .A3(new_n566_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n531_), .B1(new_n871_), .B2(KEYINPUT122), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(KEYINPUT122), .B2(new_n871_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n874_));
  INV_X1    g673(.A(G169gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  OR2_X1    g676(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n876_), .B(new_n878_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n870_), .A2(new_n475_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n842_), .A2(new_n360_), .A3(new_n633_), .A4(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n877_), .A2(new_n879_), .A3(new_n881_), .ZN(G1348gat));
  NAND3_X1  g681(.A1(new_n842_), .A2(new_n578_), .A3(new_n880_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n796_), .A2(new_n531_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n870_), .A2(new_n601_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n885_), .A2(G176gat), .A3(new_n327_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n883_), .A2(new_n359_), .B1(new_n884_), .B2(new_n886_), .ZN(G1349gat));
  AND2_X1   g686(.A1(new_n842_), .A2(new_n880_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n296_), .A2(new_n343_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n884_), .A2(new_n297_), .A3(new_n885_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n888_), .A2(new_n889_), .B1(new_n890_), .B2(new_n354_), .ZN(G1350gat));
  NAND3_X1  g690(.A1(new_n888_), .A2(new_n614_), .A3(new_n344_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n842_), .A2(new_n880_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G190gat), .B1(new_n893_), .B2(new_n267_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1351gat));
  NOR3_X1   g694(.A1(new_n587_), .A2(new_n515_), .A3(new_n479_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n848_), .B2(new_n802_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n633_), .ZN(new_n899_));
  INV_X1    g698(.A(G197gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(KEYINPUT124), .B2(new_n900_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT124), .B(G197gat), .Z(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n899_), .B2(new_n902_), .ZN(G1352gat));
  NAND2_X1  g702(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT125), .B(G204gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n898_), .A2(new_n327_), .ZN(new_n906_));
  MUX2_X1   g705(.A(new_n904_), .B(new_n905_), .S(new_n906_), .Z(G1353gat));
  AOI21_X1  g706(.A(new_n296_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n909_));
  NOR3_X1   g708(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n898_), .A2(new_n908_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n898_), .A2(new_n908_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n911_), .ZN(G1354gat));
  INV_X1    g713(.A(G218gat), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n898_), .B2(new_n624_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n263_), .A2(G218gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n898_), .A2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n917_), .A2(KEYINPUT127), .A3(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921_));
  INV_X1    g720(.A(new_n919_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n916_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n920_), .A2(new_n923_), .ZN(G1355gat));
endmodule


