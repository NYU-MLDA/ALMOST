//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n923_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_, new_n980_;
  AOI21_X1  g000(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT96), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT95), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT94), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(KEYINPUT94), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .A4(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT29), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(new_n215_), .B2(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n215_), .A2(KEYINPUT93), .A3(new_n220_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n214_), .B2(KEYINPUT1), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n221_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G141gat), .B(G148gat), .Z(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n218_), .A2(new_n219_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT28), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n213_), .A2(new_n217_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT28), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n219_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G22gat), .B(G50gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT101), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n230_), .A2(new_n219_), .ZN(new_n238_));
  OR2_X1    g037(.A1(KEYINPUT97), .A2(G197gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT97), .A2(G197gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G204gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(KEYINPUT98), .A3(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(KEYINPUT97), .A2(G197gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(KEYINPUT97), .A2(G197gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n242_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT98), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT99), .B(G204gat), .Z(new_n249_));
  OAI211_X1 g048(.A(new_n243_), .B(new_n248_), .C1(G197gat), .C2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT21), .ZN(new_n251_));
  OR2_X1    g050(.A1(KEYINPUT99), .A2(G204gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(KEYINPUT99), .A2(G204gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(G197gat), .A3(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n239_), .A2(G204gat), .A3(new_n240_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT100), .B1(new_n256_), .B2(KEYINPUT21), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT100), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT21), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n254_), .A2(new_n255_), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G211gat), .B(G218gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n251_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n256_), .A2(KEYINPUT21), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n238_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G228gat), .A2(G233gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n268_), .B(G78gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(G106gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n238_), .A2(new_n266_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n233_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n232_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n231_), .B1(new_n230_), .B2(new_n219_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT101), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n234_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n237_), .A2(new_n274_), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n278_), .B2(new_n234_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(new_n273_), .A3(new_n271_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G1gat), .B(G29gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT104), .B(KEYINPUT0), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G57gat), .B(G85gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G127gat), .B(G134gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G113gat), .B(G120gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT91), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n293_), .A2(new_n294_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT91), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n294_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n218_), .A2(new_n227_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n292_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n298_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n218_), .A2(new_n227_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n295_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n304_), .B(KEYINPUT4), .C1(new_n306_), .C2(new_n230_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n307_), .A3(KEYINPUT103), .ZN(new_n308_));
  INV_X1    g107(.A(new_n300_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n304_), .A3(new_n292_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT103), .B1(new_n302_), .B2(new_n307_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n291_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n302_), .A2(new_n307_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT103), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n316_), .A2(new_n290_), .A3(new_n310_), .A4(new_n308_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT27), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT19), .ZN(new_n322_));
  INV_X1    g121(.A(new_n265_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n264_), .B1(new_n250_), .B2(KEYINPUT21), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(new_n261_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT23), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(G183gat), .B2(G190gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G169gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT102), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(KEYINPUT102), .A3(new_n330_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G169gat), .ZN(new_n337_));
  INV_X1    g136(.A(G176gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OR3_X1    g138(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT25), .B(G183gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G190gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n344_), .A2(new_n327_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n333_), .A2(new_n334_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT20), .B1(new_n325_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n339_), .A2(new_n327_), .A3(new_n340_), .ZN(new_n348_));
  INV_X1    g147(.A(G190gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT87), .B1(new_n349_), .B2(KEYINPUT26), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT87), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G183gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT86), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G183gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n358_), .A3(KEYINPUT25), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n360_), .A2(G183gat), .B1(new_n349_), .B2(KEYINPUT26), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT88), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT88), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n354_), .A2(new_n359_), .A3(new_n364_), .A4(new_n361_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n348_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n356_), .A2(new_n358_), .A3(new_n349_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n327_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n330_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n371_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n322_), .B1(new_n347_), .B2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G8gat), .B(G36gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT18), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n378_));
  INV_X1    g177(.A(new_n371_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n266_), .B2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n322_), .B1(new_n325_), .B2(new_n346_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n373_), .A2(new_n377_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n377_), .B1(new_n373_), .B2(new_n382_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n320_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n373_), .A2(new_n382_), .A3(new_n377_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT20), .B1(new_n325_), .B2(new_n371_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n344_), .A2(new_n339_), .A3(new_n327_), .A4(new_n340_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n331_), .A2(new_n388_), .ZN(new_n389_));
  AOI211_X1 g188(.A(new_n323_), .B(new_n389_), .C1(new_n324_), .C2(new_n261_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n322_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n333_), .A2(new_n334_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n388_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n266_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n325_), .A2(new_n371_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n322_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n394_), .A2(KEYINPUT20), .A3(new_n395_), .A4(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT27), .B(new_n386_), .C1(new_n398_), .C2(new_n377_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n285_), .A2(new_n319_), .A3(new_n385_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n373_), .A2(new_n382_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n377_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT105), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n309_), .A2(new_n404_), .A3(new_n304_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n304_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT105), .B1(new_n406_), .B2(new_n300_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n292_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n290_), .B1(new_n410_), .B2(new_n307_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n403_), .A2(new_n412_), .A3(new_n386_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n317_), .A2(KEYINPUT33), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n308_), .A2(new_n310_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT33), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n290_), .A4(new_n316_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n377_), .A2(KEYINPUT32), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n391_), .B2(new_n397_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n401_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(new_n419_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n413_), .A2(new_n418_), .B1(new_n318_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n400_), .B1(new_n423_), .B2(new_n285_), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n305_), .B(KEYINPUT31), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G15gat), .B(G43gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT90), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n371_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n430_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n433_));
  INV_X1    g232(.A(G99gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n434_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n429_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n437_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n428_), .A3(new_n435_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(G71gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT92), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n443_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n426_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n446_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n448_), .A2(KEYINPUT92), .A3(new_n444_), .A4(new_n425_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n385_), .A2(new_n399_), .A3(new_n284_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT106), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n385_), .A2(new_n399_), .A3(new_n284_), .A4(KEYINPUT106), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n318_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n424_), .A2(new_n451_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G15gat), .B(G22gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G1gat), .A2(G8gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT14), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G1gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n459_), .A2(new_n460_), .A3(new_n465_), .A4(new_n461_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G29gat), .B(G36gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G43gat), .B(G50gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n471_), .A2(new_n472_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT82), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n471_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G43gat), .B(G50gat), .Z(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT82), .B1(new_n480_), .B2(new_n473_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n470_), .B1(new_n477_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n476_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(KEYINPUT82), .A3(new_n473_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n469_), .A3(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(KEYINPUT83), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n483_), .A2(new_n469_), .A3(new_n489_), .A4(new_n484_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n474_), .A2(new_n475_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n493_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n469_), .A3(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n487_), .A3(new_n482_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G113gat), .B(G141gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT84), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G169gat), .B(G197gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n491_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT85), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n491_), .A2(new_n497_), .A3(new_n504_), .A4(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n491_), .A2(new_n497_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n501_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT6), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n513_), .A2(new_n515_), .A3(KEYINPUT66), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT66), .B1(new_n513_), .B2(new_n515_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519_));
  AND2_X1   g318(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n520_));
  NOR2_X1   g319(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI22_X1  g321(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT67), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT67), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n522_), .A2(new_n526_), .A3(new_n523_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n518_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(G85gat), .ZN(new_n529_));
  INV_X1    g328(.A(G92gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G85gat), .A2(G92gat), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT8), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n528_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n513_), .A2(new_n515_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n522_), .A2(new_n537_), .A3(new_n523_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n533_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT8), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n532_), .A2(KEYINPUT9), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n542_));
  OR2_X1    g341(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n543_));
  INV_X1    g342(.A(G106gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n531_), .A2(KEYINPUT9), .A3(new_n532_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n539_), .A2(new_n540_), .B1(new_n542_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G71gat), .B(G78gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(KEYINPUT11), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n553_));
  INV_X1    g352(.A(new_n551_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n552_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n536_), .A2(new_n549_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT68), .ZN(new_n559_));
  INV_X1    g358(.A(new_n557_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT66), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n514_), .B1(G99gat), .B2(G106gat), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n512_), .A2(KEYINPUT6), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n513_), .A2(new_n515_), .A3(KEYINPUT66), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n526_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n534_), .B1(new_n568_), .B2(new_n527_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n539_), .A2(new_n540_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n548_), .A2(new_n542_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n560_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT68), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n536_), .A2(new_n574_), .A3(new_n549_), .A4(new_n557_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n559_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT64), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT69), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n536_), .A2(KEYINPUT69), .A3(new_n549_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n557_), .A2(KEYINPUT70), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT70), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n586_), .B(new_n552_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n584_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n582_), .A2(new_n583_), .A3(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n558_), .A2(new_n578_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n573_), .A2(new_n584_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G120gat), .B(G148gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n580_), .A2(new_n592_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT72), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n580_), .A2(new_n592_), .A3(KEYINPUT72), .A4(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n580_), .A2(new_n592_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n597_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n602_), .A2(KEYINPUT13), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT13), .B1(new_n602_), .B2(new_n605_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n458_), .A2(new_n511_), .A3(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT77), .B(KEYINPUT37), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT34), .Z(new_n614_));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT76), .Z(new_n617_));
  INV_X1    g416(.A(new_n492_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n536_), .A2(new_n618_), .A3(new_n549_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT75), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT75), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n536_), .A2(new_n621_), .A3(new_n618_), .A4(new_n549_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n617_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n614_), .A2(new_n615_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT73), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n582_), .A2(new_n495_), .A3(new_n494_), .A4(new_n583_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n625_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  OAI22_X1  g431(.A1(new_n628_), .A2(new_n629_), .B1(KEYINPUT36), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n629_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n632_), .B(KEYINPUT36), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(new_n627_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n612_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT17), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n585_), .A2(new_n587_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT80), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT79), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT78), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(new_n470_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n641_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n641_), .A2(new_n645_), .ZN(new_n647_));
  XOR2_X1   g446(.A(G127gat), .B(G155gat), .Z(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT16), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  OR4_X1    g450(.A1(new_n639_), .A2(new_n646_), .A3(new_n647_), .A4(new_n651_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n645_), .A2(new_n560_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n651_), .B(KEYINPUT17), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n645_), .A2(new_n560_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n633_), .A2(new_n636_), .A3(new_n612_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n638_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT81), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n610_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n463_), .A3(new_n318_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT38), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT109), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n633_), .A2(new_n636_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT107), .Z(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n458_), .B2(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n456_), .A2(new_n457_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n403_), .A2(new_n412_), .A3(new_n386_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n422_), .A2(new_n318_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n284_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n450_), .B1(new_n674_), .B2(new_n400_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT108), .B(new_n667_), .C1(new_n670_), .C2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n669_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n609_), .A2(new_n511_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n677_), .A2(new_n318_), .A3(new_n678_), .A4(new_n657_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n664_), .B1(new_n679_), .B2(G1gat), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n664_), .A3(G1gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n663_), .B1(new_n680_), .B2(new_n681_), .ZN(G1324gat));
  NAND2_X1  g481(.A1(new_n385_), .A2(new_n399_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n661_), .A2(new_n464_), .A3(new_n683_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n677_), .A2(new_n678_), .A3(new_n657_), .A4(new_n683_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(G8gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G8gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1325gat));
  INV_X1    g490(.A(G15gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n661_), .A2(new_n692_), .A3(new_n450_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n677_), .A2(new_n678_), .A3(new_n657_), .A4(new_n450_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n694_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n694_), .B2(G15gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(G1326gat));
  INV_X1    g496(.A(G22gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n661_), .A2(new_n698_), .A3(new_n285_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n677_), .A2(new_n678_), .A3(new_n657_), .A4(new_n285_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(G22gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n700_), .B2(G22gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1327gat));
  INV_X1    g503(.A(new_n666_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n657_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n610_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G29gat), .B1(new_n707_), .B2(new_n318_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n638_), .A2(KEYINPUT110), .A3(new_n658_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT110), .B1(new_n638_), .B2(new_n658_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT43), .B1(new_n458_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n658_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n637_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(KEYINPUT43), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT111), .B1(new_n458_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n718_), .B(new_n715_), .C1(new_n670_), .C2(new_n675_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n712_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n609_), .A2(new_n511_), .A3(new_n657_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(KEYINPUT44), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT44), .B1(new_n720_), .B2(new_n721_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n318_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n708_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  INV_X1    g525(.A(new_n683_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(G36gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n707_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT45), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n707_), .A2(new_n731_), .A3(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n722_), .A2(new_n723_), .A3(new_n727_), .ZN(new_n734_));
  INV_X1    g533(.A(G36gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n733_), .B(KEYINPUT46), .C1(new_n734_), .C2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1329gat));
  NAND3_X1  g539(.A1(new_n724_), .A2(G43gat), .A3(new_n450_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n707_), .A2(new_n450_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n741_), .B(new_n742_), .C1(G43gat), .C2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(G43gat), .ZN(new_n745_));
  NOR4_X1   g544(.A1(new_n722_), .A2(new_n723_), .A3(new_n745_), .A4(new_n451_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n743_), .A2(G43gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT47), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n744_), .A2(new_n748_), .ZN(G1330gat));
  AOI21_X1  g548(.A(G50gat), .B1(new_n707_), .B2(new_n285_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n285_), .A2(G50gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n724_), .B2(new_n751_), .ZN(G1331gat));
  NOR2_X1   g551(.A1(new_n608_), .A2(new_n510_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n677_), .A2(new_n657_), .A3(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G57gat), .B1(new_n754_), .B2(new_n319_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n458_), .A2(new_n510_), .A3(new_n608_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n660_), .ZN(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n318_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n759_), .ZN(G1332gat));
  INV_X1    g559(.A(G64gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n761_), .A3(new_n683_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n754_), .A2(new_n727_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G64gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G64gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(G1333gat));
  NAND3_X1  g566(.A1(new_n757_), .A2(new_n442_), .A3(new_n450_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n754_), .A2(new_n451_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G71gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G71gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1334gat));
  NOR2_X1   g572(.A1(new_n284_), .A2(G78gat), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT112), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n757_), .A2(new_n775_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n754_), .A2(new_n284_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(G78gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G78gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(G1335gat));
  NAND2_X1  g580(.A1(new_n756_), .A2(new_n706_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n529_), .A3(new_n318_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n652_), .A2(new_n656_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n753_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n720_), .A2(KEYINPUT113), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT113), .B1(new_n720_), .B2(new_n787_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n319_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n784_), .B1(new_n790_), .B2(new_n529_), .ZN(G1336gat));
  NAND3_X1  g590(.A1(new_n783_), .A2(new_n530_), .A3(new_n683_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n788_), .A2(new_n789_), .A3(new_n727_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n530_), .ZN(G1337gat));
  AND3_X1   g593(.A1(new_n720_), .A2(new_n450_), .A3(new_n787_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n450_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n796_));
  OAI22_X1  g595(.A1(new_n795_), .A2(new_n434_), .B1(new_n782_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g597(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n720_), .A2(new_n285_), .A3(new_n787_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G106gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT52), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n803_), .A3(G106gat), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n783_), .A2(new_n544_), .A3(new_n285_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n799_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n800_), .A2(new_n803_), .A3(G106gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n803_), .B1(new_n800_), .B2(G106gat), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n806_), .B(new_n799_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n807_), .A2(new_n811_), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813_));
  INV_X1    g612(.A(G113gat), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n511_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n486_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n508_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT116), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n821_), .A3(new_n508_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n496_), .A2(new_n488_), .A3(new_n482_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n506_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n589_), .A2(new_n591_), .A3(new_n559_), .A4(new_n575_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n579_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .A4(KEYINPUT55), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n592_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  AOI211_X1 g632(.A(KEYINPUT115), .B(new_n827_), .C1(new_n833_), .C2(new_n604_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n602_), .A2(new_n510_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n604_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT56), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n826_), .B1(new_n836_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n817_), .B1(new_n841_), .B2(new_n666_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n826_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n837_), .A2(new_n838_), .A3(KEYINPUT56), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n510_), .A3(new_n602_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n845_), .B2(new_n839_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n817_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n705_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n825_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n837_), .A2(KEYINPUT56), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n833_), .A2(new_n827_), .A3(new_n604_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(KEYINPUT58), .A4(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT118), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n506_), .A2(new_n824_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n851_), .A2(new_n602_), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(KEYINPUT58), .A4(new_n850_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n638_), .A2(new_n658_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n853_), .A2(new_n857_), .A3(new_n860_), .A4(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n842_), .A2(new_n848_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n785_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n607_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n602_), .A2(KEYINPUT13), .A3(new_n605_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n511_), .A3(new_n866_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n867_), .A2(new_n659_), .A3(KEYINPUT54), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n606_), .A2(new_n607_), .A3(new_n510_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n713_), .A2(new_n785_), .A3(new_n637_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n868_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n864_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n456_), .A2(new_n318_), .A3(new_n450_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(KEYINPUT120), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n873_), .B1(new_n863_), .B2(new_n785_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n876_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n816_), .B1(new_n880_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n881_), .A2(new_n511_), .A3(new_n876_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(G113gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n875_), .A2(new_n510_), .A3(new_n877_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(KEYINPUT119), .A3(new_n814_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n813_), .B1(new_n884_), .B2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT59), .B1(new_n882_), .B2(KEYINPUT120), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893_));
  NOR4_X1   g692(.A1(new_n881_), .A2(new_n893_), .A3(new_n879_), .A4(new_n876_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n815_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n895_), .A2(KEYINPUT121), .A3(new_n887_), .A4(new_n889_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n891_), .A2(new_n896_), .ZN(G1340gat));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n608_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n882_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n608_), .B1(new_n880_), .B2(new_n883_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n898_), .ZN(G1341gat));
  NAND2_X1  g701(.A1(new_n880_), .A2(new_n883_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(G127gat), .A3(new_n657_), .ZN(new_n904_));
  INV_X1    g703(.A(G127gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n875_), .A2(new_n877_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n785_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n907_), .A2(KEYINPUT122), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(KEYINPUT122), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n904_), .A2(new_n908_), .A3(new_n909_), .ZN(G1342gat));
  INV_X1    g709(.A(G134gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(new_n906_), .B2(new_n667_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT123), .B(new_n911_), .C1(new_n906_), .C2(new_n667_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n714_), .A2(new_n911_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n903_), .B2(new_n917_), .ZN(G1343gat));
  NAND3_X1  g717(.A1(new_n727_), .A2(new_n318_), .A3(new_n285_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n881_), .A2(new_n450_), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n510_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n609_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g723(.A1(new_n920_), .A2(new_n657_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT61), .B(G155gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1346gat));
  AOI21_X1  g726(.A(G162gat), .B1(new_n920_), .B2(new_n668_), .ZN(new_n928_));
  INV_X1    g727(.A(G162gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n711_), .A2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n920_), .B2(new_n930_), .ZN(G1347gat));
  NAND2_X1  g730(.A1(new_n875_), .A2(new_n683_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n457_), .A2(new_n284_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n510_), .ZN(new_n935_));
  OAI211_X1 g734(.A(KEYINPUT62), .B(G169gat), .C1(new_n935_), .C2(KEYINPUT22), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n881_), .A2(new_n727_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n933_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n511_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT22), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n937_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n337_), .B1(new_n941_), .B2(new_n937_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n936_), .B1(new_n943_), .B2(new_n944_), .ZN(G1348gat));
  NOR2_X1   g744(.A1(new_n940_), .A2(new_n608_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n338_), .ZN(G1349gat));
  INV_X1    g746(.A(new_n342_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n938_), .A2(new_n657_), .A3(new_n948_), .A4(new_n939_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n932_), .A2(new_n785_), .A3(new_n933_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n356_), .A2(new_n358_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n949_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(KEYINPUT124), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954_));
  OAI211_X1 g753(.A(new_n954_), .B(new_n949_), .C1(new_n950_), .C2(new_n951_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n955_), .ZN(G1350gat));
  NAND3_X1  g755(.A1(new_n934_), .A2(new_n343_), .A3(new_n668_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n938_), .A2(new_n861_), .A3(new_n939_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959_));
  AND3_X1   g758(.A1(new_n958_), .A2(new_n959_), .A3(G190gat), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n959_), .B1(new_n958_), .B2(G190gat), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n957_), .B1(new_n960_), .B2(new_n961_), .ZN(G1351gat));
  NOR3_X1   g761(.A1(new_n450_), .A2(new_n318_), .A3(new_n284_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n938_), .A2(new_n963_), .ZN(new_n964_));
  INV_X1    g763(.A(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(new_n510_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g766(.A1(new_n964_), .A2(new_n608_), .ZN(new_n968_));
  MUX2_X1   g767(.A(G204gat), .B(new_n249_), .S(new_n968_), .Z(G1353gat));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970_));
  INV_X1    g769(.A(G211gat), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n657_), .B1(new_n970_), .B2(new_n971_), .ZN(new_n972_));
  XOR2_X1   g771(.A(new_n972_), .B(KEYINPUT126), .Z(new_n973_));
  NAND2_X1  g772(.A1(new_n965_), .A2(new_n973_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n970_), .A2(new_n971_), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n974_), .B(new_n975_), .ZN(G1354gat));
  AND3_X1   g775(.A1(new_n965_), .A2(G218gat), .A3(new_n861_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n964_), .A2(new_n667_), .ZN(new_n978_));
  OR2_X1    g777(.A1(new_n978_), .A2(KEYINPUT127), .ZN(new_n979_));
  AOI21_X1  g778(.A(G218gat), .B1(new_n978_), .B2(KEYINPUT127), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n977_), .B1(new_n979_), .B2(new_n980_), .ZN(G1355gat));
endmodule


