//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n970_, new_n971_,
    new_n972_, new_n974_, new_n975_, new_n976_, new_n978_, new_n979_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n986_, new_n988_,
    new_n989_, new_n990_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  AND2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT88), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n208_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n205_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n204_), .B1(new_n202_), .B2(KEYINPUT1), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n222_), .A2(new_n223_), .B1(G141gat), .B2(G148gat), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n220_), .A2(new_n224_), .A3(KEYINPUT87), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT87), .B1(new_n220_), .B2(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n217_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT89), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n217_), .B(new_n229_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n228_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n220_), .A2(new_n224_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n220_), .A2(new_n224_), .A3(KEYINPUT87), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n215_), .A2(new_n216_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n238_), .A2(new_n239_), .B1(new_n240_), .B2(new_n205_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n233_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n235_), .A2(KEYINPUT4), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n228_), .A2(new_n230_), .A3(new_n234_), .A4(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n243_), .A2(KEYINPUT97), .A3(new_n245_), .A4(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n235_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n245_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT97), .B1(new_n252_), .B2(new_n243_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT103), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT98), .B(KEYINPUT0), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT99), .ZN(new_n257_));
  XOR2_X1   g056(.A(G1gat), .B(G29gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G57gat), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n254_), .A2(new_n255_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT97), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n235_), .A2(KEYINPUT4), .A3(new_n242_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(new_n251_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n266_), .A2(new_n262_), .A3(new_n249_), .A4(new_n248_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT103), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n261_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT102), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT22), .B(G169gat), .ZN(new_n272_));
  INV_X1    g071(.A(G176gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n278_));
  INV_X1    g077(.A(G183gat), .ZN(new_n279_));
  INV_X1    g078(.A(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n278_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n274_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285_));
  INV_X1    g084(.A(G169gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(new_n273_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT26), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n280_), .A2(KEYINPUT26), .ZN(new_n291_));
  AND2_X1   g090(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n290_), .B(new_n291_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n286_), .A2(new_n273_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(KEYINPUT24), .A3(new_n283_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT95), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n288_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(KEYINPUT95), .A3(new_n296_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n284_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G218gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G211gat), .ZN(new_n303_));
  INV_X1    g102(.A(G211gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G218gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT90), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT90), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n303_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G197gat), .A2(G204gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G197gat), .A2(G204gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(KEYINPUT21), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT21), .ZN(new_n314_));
  INV_X1    g113(.A(new_n312_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(new_n310_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n307_), .A2(new_n309_), .A3(new_n313_), .A4(new_n316_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n315_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n303_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n308_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT92), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT92), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n317_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n301_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(KEYINPUT91), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT81), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n288_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n287_), .A2(new_n277_), .A3(KEYINPUT81), .A4(new_n278_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT25), .B1(new_n279_), .B2(KEYINPUT79), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(G183gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n332_), .B(new_n335_), .C1(new_n336_), .C2(new_n291_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n289_), .A2(G190gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n290_), .B1(new_n338_), .B2(KEYINPUT80), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n296_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(KEYINPUT82), .A2(G169gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(KEYINPUT82), .A2(G169gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT83), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n277_), .A2(new_n281_), .A3(new_n347_), .A4(new_n278_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n341_), .A2(new_n344_), .A3(new_n342_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n282_), .A2(KEYINPUT83), .ZN(new_n351_));
  OAI22_X1  g150(.A1(new_n331_), .A2(new_n340_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT91), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n317_), .A2(new_n321_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n327_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n326_), .A2(new_n355_), .A3(KEYINPUT20), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT19), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n352_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n354_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n353_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n322_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n301_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n358_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n363_), .A2(new_n365_), .A3(KEYINPUT20), .A4(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n271_), .B1(new_n359_), .B2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT102), .B1(new_n356_), .B2(new_n358_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n358_), .B1(new_n301_), .B2(new_n364_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(KEYINPUT20), .A3(new_n355_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n352_), .B1(new_n354_), .B2(new_n327_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n301_), .A2(new_n364_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n372_), .B1(new_n376_), .B2(new_n366_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n382_));
  MUX2_X1   g181(.A(new_n370_), .B(new_n377_), .S(new_n382_), .Z(new_n383_));
  INV_X1    g182(.A(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n377_), .A2(new_n384_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n381_), .B(new_n372_), .C1(new_n376_), .C2(new_n366_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n235_), .A2(KEYINPUT101), .A3(new_n242_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT101), .B1(new_n235_), .B2(new_n242_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n244_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n247_), .A2(new_n244_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n261_), .B1(new_n265_), .B2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n385_), .B(new_n386_), .C1(new_n389_), .C2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT100), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n267_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n394_), .B2(KEYINPUT33), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n267_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n270_), .A2(new_n383_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT93), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n228_), .A2(KEYINPUT29), .A3(new_n230_), .ZN(new_n400_));
  AND2_X1   g199(.A1(G228gat), .A2(G233gat), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n361_), .A2(new_n401_), .A3(new_n362_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n317_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n324_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n405_));
  OAI22_X1  g204(.A1(new_n241_), .A2(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n400_), .A2(new_n402_), .B1(new_n406_), .B2(new_n401_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n399_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT29), .B1(new_n228_), .B2(new_n230_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G22gat), .B(G50gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n412_), .B(KEYINPUT28), .Z(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n411_), .B(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT94), .B1(new_n410_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n400_), .A2(new_n402_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n406_), .A2(new_n401_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n409_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT93), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n411_), .B(new_n413_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT94), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n416_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n407_), .B(new_n408_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n416_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n384_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT104), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT104), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n432_), .B(new_n384_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n386_), .A2(KEYINPUT27), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT105), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n385_), .A2(new_n386_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT27), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT105), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n431_), .A2(new_n441_), .A3(new_n433_), .A4(new_n435_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n437_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n269_), .B1(KEYINPUT103), .B2(new_n267_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n267_), .A2(KEYINPUT103), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n429_), .ZN(new_n447_));
  OAI22_X1  g246(.A1(new_n398_), .A2(new_n429_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT31), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT84), .B1(new_n233_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(new_n449_), .B2(new_n233_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(G43gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n451_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455_));
  INV_X1    g254(.A(G15gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT30), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n454_), .B(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n352_), .B(KEYINPUT85), .Z(new_n461_));
  OR2_X1    g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n461_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n416_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n425_), .B1(new_n416_), .B2(new_n423_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n437_), .A2(new_n467_), .A3(new_n440_), .A4(new_n442_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n446_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT106), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n442_), .A2(new_n440_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n434_), .B1(new_n430_), .B2(KEYINPUT104), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n441_), .B1(new_n473_), .B2(new_n433_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT106), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n270_), .A2(new_n464_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n467_), .A4(new_n477_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n448_), .A2(new_n464_), .B1(new_n471_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G230gat), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT64), .ZN(new_n482_));
  INV_X1    g281(.A(G99gat), .ZN(new_n483_));
  INV_X1    g282(.A(G106gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT7), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT6), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n482_), .A2(new_n492_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n486_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT66), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT8), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT65), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n496_), .A2(KEYINPUT65), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499_));
  INV_X1    g298(.A(G85gat), .ZN(new_n500_));
  INV_X1    g299(.A(G92gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n498_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n494_), .A2(new_n497_), .A3(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n484_), .A3(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n502_), .A2(KEYINPUT9), .A3(new_n499_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n499_), .A2(KEYINPUT9), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n491_), .A2(new_n507_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n497_), .B1(new_n494_), .B2(new_n503_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT67), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G57gat), .B(G64gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT11), .ZN(new_n516_));
  XOR2_X1   g315(.A(G71gat), .B(G78gat), .Z(new_n517_));
  INV_X1    g316(.A(G64gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G57gat), .ZN(new_n519_));
  INV_X1    g318(.A(G57gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G64gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n521_), .A3(KEYINPUT11), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n514_), .A2(KEYINPUT11), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n516_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n494_), .A2(new_n503_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n497_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n510_), .A4(new_n504_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n513_), .A2(new_n525_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n525_), .B1(new_n513_), .B2(new_n530_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n481_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G120gat), .B(G148gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT5), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(KEYINPUT12), .B(new_n516_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n541_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT68), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n544_), .B(new_n541_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n546_), .B(new_n531_), .C1(KEYINPUT12), .C2(new_n533_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n534_), .B(new_n539_), .C1(new_n547_), .C2(new_n481_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n513_), .A2(new_n530_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n551_), .A2(new_n525_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n513_), .A2(new_n530_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n525_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(new_n557_), .A3(new_n480_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n558_), .A2(KEYINPUT69), .A3(new_n534_), .A4(new_n539_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n550_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n534_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n538_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n560_), .A2(KEYINPUT13), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT13), .B1(new_n560_), .B2(new_n562_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G29gat), .B(G36gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G43gat), .B(G50gat), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G43gat), .B(G50gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n570_), .A2(KEYINPUT15), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT15), .B1(new_n570_), .B2(new_n572_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(G22gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n456_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G15gat), .A2(G22gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G1gat), .A2(G8gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT14), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n585_));
  INV_X1    g384(.A(G1gat), .ZN(new_n586_));
  INV_X1    g385(.A(G8gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n585_), .B1(new_n588_), .B2(new_n582_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n585_), .A3(new_n582_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n584_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n579_), .A2(new_n580_), .B1(KEYINPUT14), .B2(new_n582_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n589_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n577_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n593_), .B2(new_n589_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n591_), .A3(new_n584_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n576_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n575_), .A2(new_n596_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n570_), .A2(new_n572_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n576_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n576_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n601_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT78), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n600_), .A2(new_n604_), .A3(new_n605_), .A4(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n600_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT78), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n596_), .A2(new_n599_), .A3(new_n572_), .A4(new_n570_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n606_), .B1(new_n604_), .B2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G169gat), .B(G197gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n607_), .B(new_n617_), .C1(new_n609_), .C2(new_n611_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n566_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n479_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT34), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(KEYINPUT35), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n528_), .A2(new_n510_), .A3(new_n504_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n575_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n628_), .B2(KEYINPUT71), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT71), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n627_), .A2(new_n575_), .A3(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n513_), .A2(new_n530_), .A3(new_n601_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT72), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n513_), .A2(new_n530_), .A3(KEYINPUT72), .A4(new_n601_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n625_), .A2(KEYINPUT35), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT70), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT36), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G190gat), .B(G218gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT73), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G134gat), .B(G162gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n626_), .B(new_n641_), .C1(new_n627_), .C2(new_n575_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n637_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n642_), .A2(new_n643_), .A3(new_n647_), .A4(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n643_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n647_), .A2(new_n643_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n640_), .B1(new_n632_), .B2(new_n637_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n649_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n651_), .B(new_n652_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT37), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n650_), .A2(new_n655_), .A3(KEYINPUT37), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n596_), .A2(new_n599_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(G231gat), .A2(G233gat), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n525_), .B(new_n663_), .Z(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n525_), .B(new_n663_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n661_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(G127gat), .B(G155gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(G183gat), .B(G211gat), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n672_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(KEYINPUT17), .A3(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n668_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n674_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT17), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n675_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n676_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n660_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n623_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n586_), .A3(new_n270_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT38), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n656_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n479_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n622_), .A2(new_n683_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G1gat), .B1(new_n693_), .B2(new_n446_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n687_), .A2(new_n688_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n689_), .A2(new_n694_), .A3(new_n695_), .ZN(G1324gat));
  NAND3_X1  g495(.A1(new_n686_), .A2(new_n587_), .A3(new_n443_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n693_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n443_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT39), .ZN(new_n700_));
  OAI21_X1  g499(.A(G8gat), .B1(new_n700_), .B2(KEYINPUT107), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n699_), .A2(new_n702_), .B1(KEYINPUT107), .B2(new_n700_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(KEYINPUT107), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n704_), .B(new_n701_), .C1(new_n698_), .C2(new_n443_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n697_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT40), .B(new_n697_), .C1(new_n703_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1325gat));
  NAND3_X1  g509(.A1(new_n686_), .A2(new_n456_), .A3(new_n469_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G15gat), .B1(new_n693_), .B2(new_n464_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(new_n713_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT108), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n718_), .B(new_n711_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1326gat));
  OAI21_X1  g519(.A(G22gat), .B1(new_n693_), .B2(new_n467_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT42), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n686_), .A2(new_n578_), .A3(new_n429_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1327gat));
  NOR2_X1   g523(.A1(new_n656_), .A2(new_n682_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n623_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G29gat), .B1(new_n726_), .B2(new_n270_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n659_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT37), .B1(new_n650_), .B2(new_n655_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT43), .B1(new_n479_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n471_), .A2(new_n478_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n443_), .A2(new_n447_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n270_), .A2(new_n383_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n395_), .A2(new_n397_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n429_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n464_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n732_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n739_), .A3(new_n660_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n731_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n621_), .A2(new_n683_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT44), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n745_), .B(new_n742_), .C1(new_n731_), .C2(new_n740_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n270_), .A2(G29gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n727_), .B1(new_n747_), .B2(new_n748_), .ZN(G1328gat));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n750_));
  INV_X1    g549(.A(G36gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n747_), .B2(new_n443_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n623_), .A2(new_n751_), .A3(new_n443_), .A4(new_n725_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n752_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n755_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n744_), .A2(new_n746_), .A3(new_n475_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n757_), .B(KEYINPUT46), .C1(new_n758_), .C2(new_n751_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(G1329gat));
  INV_X1    g559(.A(G43gat), .ZN(new_n761_));
  NOR4_X1   g560(.A1(new_n744_), .A2(new_n746_), .A3(new_n761_), .A4(new_n464_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G43gat), .B1(new_n726_), .B2(new_n469_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT47), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n464_), .A2(new_n761_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n747_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n764_), .A2(new_n768_), .ZN(G1330gat));
  AOI21_X1  g568(.A(G50gat), .B1(new_n726_), .B2(new_n429_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n429_), .A2(G50gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n747_), .B2(new_n771_), .ZN(G1331gat));
  NAND3_X1  g571(.A1(new_n616_), .A2(new_n682_), .A3(new_n618_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n565_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n691_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(G57gat), .A3(new_n270_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n777_), .A2(new_n778_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n479_), .A2(new_n619_), .A3(new_n565_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n684_), .ZN(new_n782_));
  AOI21_X1  g581(.A(G57gat), .B1(new_n782_), .B2(new_n270_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n779_), .A2(new_n780_), .A3(new_n783_), .ZN(G1332gat));
  NAND2_X1  g583(.A1(new_n443_), .A2(new_n518_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT111), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G64gat), .B1(new_n775_), .B2(new_n475_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(KEYINPUT48), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(KEYINPUT48), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT112), .B(new_n787_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1333gat));
  INV_X1    g594(.A(G71gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n782_), .A2(new_n796_), .A3(new_n469_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n776_), .B2(new_n469_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n799_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(G1334gat));
  OAI21_X1  g601(.A(G78gat), .B1(new_n775_), .B2(new_n467_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(G78gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n782_), .A2(new_n806_), .A3(new_n429_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1335gat));
  NOR3_X1   g607(.A1(new_n565_), .A2(new_n682_), .A3(new_n619_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n741_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(G85gat), .B1(new_n810_), .B2(new_n446_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n781_), .A2(new_n725_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n270_), .A2(new_n500_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(G1336gat));
  OAI21_X1  g615(.A(G92gat), .B1(new_n810_), .B2(new_n475_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n443_), .A2(new_n501_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n814_), .B2(new_n818_), .ZN(G1337gat));
  NAND3_X1  g618(.A1(new_n469_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n814_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n810_), .A2(new_n464_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(new_n483_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT51), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n825_));
  OAI221_X1 g624(.A(new_n825_), .B1(new_n822_), .B2(new_n483_), .C1(new_n814_), .C2(new_n820_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1338gat));
  NAND3_X1  g626(.A1(new_n741_), .A2(new_n429_), .A3(new_n809_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n484_), .B1(new_n829_), .B2(KEYINPUT52), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(KEYINPUT52), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n828_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n429_), .A2(new_n484_), .ZN(new_n834_));
  OAI22_X1  g633(.A1(new_n832_), .A2(new_n833_), .B1(new_n814_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT53), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837_));
  OAI221_X1 g636(.A(new_n837_), .B1(new_n814_), .B2(new_n834_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1339gat));
  NAND2_X1  g638(.A1(new_n560_), .A2(new_n562_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT13), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n773_), .B(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n560_), .A2(KEYINPUT13), .A3(new_n562_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n842_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n846_), .B2(new_n660_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n565_), .A2(new_n730_), .A3(new_n848_), .A4(new_n844_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n560_), .A2(new_n619_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n545_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n544_), .B1(new_n627_), .B2(new_n541_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n531_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT12), .B1(new_n553_), .B2(new_n554_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n481_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n547_), .A2(new_n481_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(KEYINPUT55), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n547_), .A2(new_n859_), .A3(new_n481_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n538_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT56), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n480_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n558_), .B1(new_n864_), .B2(new_n859_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n857_), .A2(new_n856_), .A3(KEYINPUT55), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT56), .A3(new_n538_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n851_), .B1(new_n863_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n606_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n604_), .B2(new_n610_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n872_));
  OR3_X1    g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n615_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n600_), .A2(new_n604_), .A3(new_n870_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n871_), .B2(new_n615_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n616_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n656_), .B1(new_n869_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(KEYINPUT57), .B(new_n656_), .C1(new_n869_), .C2(new_n878_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n877_), .B1(new_n550_), .B2(new_n559_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT56), .B1(new_n867_), .B2(new_n538_), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n862_), .B(new_n539_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT58), .B(new_n883_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n660_), .A3(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n881_), .A2(new_n882_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n850_), .B1(new_n891_), .B2(new_n683_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n468_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n446_), .A2(new_n464_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n892_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(G113gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n619_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n896_), .A2(KEYINPUT59), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(KEYINPUT59), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n620_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n898_), .B1(new_n901_), .B2(new_n897_), .ZN(G1340gat));
  OR2_X1    g701(.A1(new_n565_), .A2(KEYINPUT60), .ZN(new_n903_));
  INV_X1    g702(.A(G120gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n896_), .B(new_n905_), .C1(KEYINPUT60), .C2(new_n904_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n565_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT119), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n906_), .B(new_n910_), .C1(new_n907_), .C2(new_n904_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1341gat));
  AOI21_X1  g711(.A(G127gat), .B1(new_n896_), .B2(new_n682_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n913_), .A2(KEYINPUT120), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(KEYINPUT120), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n899_), .A2(new_n900_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n682_), .A2(G127gat), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n914_), .A2(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(G1342gat));
  INV_X1    g717(.A(G134gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n896_), .A2(new_n919_), .A3(new_n690_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n730_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n919_), .ZN(G1343gat));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n620_), .B1(new_n550_), .B2(new_n559_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n878_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n690_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n889_), .A2(new_n660_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n863_), .A2(new_n868_), .ZN(new_n929_));
  AOI21_X1  g728(.A(KEYINPUT58), .B1(new_n929_), .B2(new_n883_), .ZN(new_n930_));
  OAI22_X1  g729(.A1(new_n927_), .A2(KEYINPUT57), .B1(new_n928_), .B2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n882_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n683_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n850_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n469_), .B1(new_n933_), .B2(new_n934_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n475_), .A2(new_n429_), .A3(new_n270_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n923_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n938_));
  NOR4_X1   g737(.A1(new_n892_), .A2(KEYINPUT121), .A3(new_n469_), .A4(new_n936_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n620_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n211_), .ZN(G1344gat));
  NOR2_X1   g741(.A1(new_n940_), .A2(new_n565_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(new_n212_), .ZN(G1345gat));
  OAI21_X1  g743(.A(new_n682_), .B1(new_n938_), .B2(new_n939_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(KEYINPUT122), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n947_), .B(new_n682_), .C1(new_n938_), .C2(new_n939_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(KEYINPUT61), .B(G155gat), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n946_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n946_), .B2(new_n948_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1346gat));
  OAI21_X1  g751(.A(G162gat), .B1(new_n940_), .B2(new_n730_), .ZN(new_n953_));
  OR2_X1    g752(.A1(new_n656_), .A2(G162gat), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n940_), .B2(new_n954_), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n475_), .A2(new_n470_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(KEYINPUT123), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n892_), .A2(new_n429_), .A3(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n619_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n959_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n960_));
  INV_X1    g759(.A(new_n272_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n961_), .B2(new_n959_), .ZN(new_n962_));
  AOI21_X1  g761(.A(KEYINPUT62), .B1(new_n959_), .B2(G169gat), .ZN(new_n963_));
  OR2_X1    g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1348gat));
  INV_X1    g763(.A(new_n958_), .ZN(new_n965_));
  AOI211_X1 g764(.A(new_n565_), .B(new_n965_), .C1(KEYINPUT124), .C2(new_n273_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(KEYINPUT124), .B(G176gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n967_), .B1(new_n958_), .B2(new_n566_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n966_), .A2(new_n968_), .ZN(G1349gat));
  NAND2_X1  g768(.A1(new_n958_), .A2(new_n682_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(G183gat), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n292_), .A2(new_n293_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n970_), .B2(new_n972_), .ZN(G1350gat));
  OAI21_X1  g772(.A(G190gat), .B1(new_n965_), .B2(new_n730_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n690_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n975_), .B(KEYINPUT125), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n974_), .B1(new_n965_), .B2(new_n976_), .ZN(G1351gat));
  NOR4_X1   g776(.A1(new_n892_), .A2(new_n447_), .A3(new_n475_), .A4(new_n469_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n978_), .A2(new_n619_), .ZN(new_n979_));
  XNOR2_X1  g778(.A(new_n979_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g779(.A1(new_n978_), .A2(new_n566_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g781(.A(new_n683_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n983_));
  XOR2_X1   g782(.A(new_n983_), .B(KEYINPUT126), .Z(new_n984_));
  NAND2_X1  g783(.A1(new_n978_), .A2(new_n984_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n986_));
  XOR2_X1   g785(.A(new_n985_), .B(new_n986_), .Z(G1354gat));
  NAND3_X1  g786(.A1(new_n978_), .A2(new_n302_), .A3(new_n690_), .ZN(new_n988_));
  AND2_X1   g787(.A1(new_n978_), .A2(new_n660_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n988_), .B1(new_n989_), .B2(new_n302_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n990_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


