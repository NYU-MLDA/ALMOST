//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n849_, new_n850_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_;
  INV_X1    g000(.A(G85gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT67), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  INV_X1    g016(.A(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT7), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(KEYINPUT65), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT65), .B1(new_n224_), .B2(new_n217_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n222_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n206_), .B1(new_n216_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n212_), .A2(new_n213_), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n222_), .B(new_n230_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n206_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n204_), .A2(KEYINPUT9), .A3(new_n205_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n230_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT10), .B(G99gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(G106gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n234_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n235_), .A2(new_n236_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n219_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n241_), .A2(new_n243_), .A3(KEYINPUT64), .A4(new_n230_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n229_), .A2(new_n233_), .B1(new_n240_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G57gat), .ZN(new_n246_));
  INV_X1    g045(.A(G64gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G57gat), .A2(G64gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G71gat), .A2(G78gat), .ZN(new_n252_));
  INV_X1    g051(.A(G71gat), .ZN(new_n253_));
  INV_X1    g052(.A(G78gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT68), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n249_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n251_), .A2(new_n259_), .A3(new_n252_), .A4(new_n255_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n257_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n258_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n245_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n244_), .A2(new_n240_), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n266_));
  NOR3_X1   g065(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n267_));
  OAI22_X1  g066(.A1(new_n266_), .A2(new_n223_), .B1(new_n267_), .B2(KEYINPUT65), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n211_), .A2(new_n268_), .A3(new_n222_), .A4(new_n215_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n232_), .B1(new_n269_), .B2(new_n206_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n231_), .A2(new_n232_), .A3(new_n206_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n265_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n261_), .A2(new_n262_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n264_), .A2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(G230gat), .A2(G233gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n272_), .A2(KEYINPUT12), .A3(new_n273_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT12), .B1(new_n272_), .B2(new_n273_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n276_), .B1(new_n245_), .B2(new_n263_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n278_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT12), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n274_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n272_), .A2(KEYINPUT12), .A3(new_n273_), .ZN(new_n286_));
  AND4_X1   g085(.A1(new_n278_), .A2(new_n285_), .A3(new_n282_), .A4(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n277_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G120gat), .B(G148gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(G176gat), .B(G204gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n295_));
  INV_X1    g094(.A(new_n293_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n277_), .B(new_n296_), .C1(new_n283_), .C2(new_n287_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n288_), .A2(KEYINPUT71), .A3(new_n293_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT13), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G29gat), .B(G36gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G43gat), .B(G50gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G15gat), .B(G22gat), .ZN(new_n310_));
  INV_X1    g109(.A(G1gat), .ZN(new_n311_));
  INV_X1    g110(.A(G8gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT14), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G8gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n309_), .B(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(G229gat), .A2(G233gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n309_), .A2(KEYINPUT15), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT15), .ZN(new_n322_));
  INV_X1    g121(.A(new_n308_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n307_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n307_), .A2(new_n323_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n322_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  MUX2_X1   g126(.A(new_n309_), .B(new_n327_), .S(new_n316_), .Z(new_n328_));
  OAI21_X1  g127(.A(new_n320_), .B1(new_n328_), .B2(new_n319_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G113gat), .B(G141gat), .ZN(new_n330_));
  INV_X1    g129(.A(G169gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G197gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT79), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n329_), .B(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n304_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT37), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n327_), .A2(new_n272_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G232gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT34), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n245_), .A2(new_n309_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n340_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n343_), .A2(new_n345_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n349_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n340_), .A2(new_n351_), .A3(new_n346_), .A4(new_n347_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n350_), .A2(KEYINPUT76), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT76), .B1(new_n350_), .B2(new_n352_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G190gat), .B(G218gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G134gat), .ZN(new_n356_));
  INV_X1    g155(.A(G162gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT36), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n353_), .A2(new_n354_), .A3(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n350_), .A2(new_n352_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n358_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(KEYINPUT36), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n339_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n364_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n367_), .B(KEYINPUT37), .C1(new_n362_), .C2(new_n360_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n273_), .B(new_n317_), .ZN(new_n371_));
  AND2_X1   g170(.A1(G231gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n373_), .A2(KEYINPUT77), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT16), .B(G183gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G211gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G127gat), .B(G155gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  OR3_X1    g177(.A1(new_n374_), .A2(KEYINPUT17), .A3(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n374_), .A2(new_n378_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n373_), .A2(new_n378_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT17), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n379_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n370_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT78), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT98), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388_));
  OR3_X1    g187(.A1(new_n388_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT81), .B1(new_n388_), .B2(KEYINPUT23), .ZN(new_n390_));
  INV_X1    g189(.A(new_n388_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT80), .B(KEYINPUT23), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n389_), .B(new_n390_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(G183gat), .B2(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT22), .B(G169gat), .ZN(new_n397_));
  INV_X1    g196(.A(G176gat), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n388_), .A2(KEYINPUT23), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n405_), .B2(new_n395_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT25), .B(G183gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT26), .B(G190gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n400_), .B1(new_n402_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G197gat), .B(G204gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT89), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT21), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G211gat), .B(G218gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n415_), .B2(KEYINPUT89), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n418_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n412_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT91), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n424_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n410_), .A2(new_n393_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(G183gat), .A2(G190gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n399_), .B1(new_n402_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n427_), .A2(KEYINPUT20), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G226gat), .A2(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT19), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G8gat), .B(G36gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n428_), .A2(new_n433_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT20), .B1(new_n412_), .B2(new_n424_), .ZN(new_n446_));
  OR3_X1    g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n437_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n438_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n444_), .B1(new_n438_), .B2(new_n447_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n387_), .B1(new_n450_), .B2(KEYINPUT27), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n438_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n437_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n443_), .B(KEYINPUT96), .Z(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n438_), .A2(KEYINPUT97), .A3(new_n444_), .A4(new_n447_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n454_), .A2(KEYINPUT27), .A3(new_n458_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT27), .ZN(new_n461_));
  OAI211_X1 g260(.A(KEYINPUT98), .B(new_n461_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n451_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(G155gat), .A2(G162gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT1), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G141gat), .ZN(new_n469_));
  INV_X1    g268(.A(G148gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n464_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT85), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n466_), .B(KEYINPUT86), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n471_), .A2(KEYINPUT3), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(KEYINPUT3), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT2), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n476_), .A2(new_n477_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n474_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G127gat), .B(G134gat), .ZN(new_n484_));
  INV_X1    g283(.A(G113gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G120gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n483_), .B(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G225gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT94), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(KEYINPUT4), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(KEYINPUT93), .ZN(new_n494_));
  INV_X1    g293(.A(new_n483_), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n495_), .A2(KEYINPUT4), .A3(new_n488_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(KEYINPUT93), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n492_), .B1(new_n498_), .B2(new_n491_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT0), .B(G57gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(G85gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(G1gat), .B(G29gat), .Z(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  NOR2_X1   g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n503_), .ZN(new_n505_));
  AOI211_X1 g304(.A(new_n505_), .B(new_n492_), .C1(new_n498_), .C2(new_n491_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G22gat), .B(G50gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT87), .B1(new_n483_), .B2(KEYINPUT29), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n483_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n510_), .A2(G228gat), .A3(G233gat), .A4(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n483_), .A2(new_n511_), .A3(KEYINPUT29), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n428_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n510_), .A2(new_n424_), .B1(G228gat), .B2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT28), .B(G78gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n515_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n483_), .A2(KEYINPUT29), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G106gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n518_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n521_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n509_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n432_), .B(KEYINPUT30), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G227gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G15gat), .B(G43gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT82), .ZN(new_n531_));
  XOR2_X1   g330(.A(G71gat), .B(G99gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n529_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT84), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n488_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(KEYINPUT84), .A3(new_n535_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n536_), .A2(new_n537_), .A3(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n519_), .A2(new_n522_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n521_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n508_), .A3(new_n523_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n526_), .A2(new_n545_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n545_), .B1(new_n526_), .B2(new_n549_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n463_), .B(new_n507_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n499_), .B2(new_n503_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT33), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT95), .ZN(new_n556_));
  INV_X1    g355(.A(new_n491_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n497_), .A2(new_n496_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(new_n494_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n505_), .B(new_n556_), .C1(new_n559_), .C2(new_n492_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n489_), .A2(new_n491_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n503_), .B(new_n561_), .C1(new_n498_), .C2(new_n491_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n554_), .A2(new_n560_), .A3(new_n450_), .A4(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n444_), .A2(KEYINPUT32), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n438_), .A2(new_n447_), .A3(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n456_), .A2(KEYINPUT32), .A3(new_n444_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n565_), .B(new_n566_), .C1(new_n504_), .C2(new_n506_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n526_), .A2(new_n549_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n545_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n552_), .A2(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n338_), .A2(new_n386_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n507_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n311_), .A3(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT100), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n338_), .A2(new_n571_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n353_), .A2(new_n354_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n367_), .B1(new_n581_), .B2(new_n360_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n383_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G1gat), .B1(new_n585_), .B2(new_n507_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n578_), .B(new_n586_), .C1(new_n576_), .C2(new_n574_), .ZN(G1324gat));
  INV_X1    g386(.A(KEYINPUT40), .ZN(new_n588_));
  INV_X1    g387(.A(new_n463_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n580_), .A2(new_n589_), .A3(new_n584_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(G8gat), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT39), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n572_), .A2(new_n312_), .A3(new_n589_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT101), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n588_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n596_), .B(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n600_), .A2(KEYINPUT40), .A3(new_n594_), .A4(new_n593_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(G1325gat));
  INV_X1    g401(.A(G15gat), .ZN(new_n603_));
  INV_X1    g402(.A(new_n545_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n572_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G15gat), .B1(new_n585_), .B2(new_n545_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT41), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(G1326gat));
  OAI21_X1  g409(.A(G22gat), .B1(new_n585_), .B2(new_n569_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT102), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT102), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n613_), .B(G22gat), .C1(new_n585_), .C2(new_n569_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT42), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(KEYINPUT42), .A3(new_n614_), .ZN(new_n618_));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n569_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n572_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(new_n618_), .A3(new_n621_), .ZN(G1327gat));
  NOR2_X1   g421(.A1(new_n384_), .A2(new_n582_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n579_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(G29gat), .B1(new_n625_), .B2(new_n573_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n571_), .A2(new_n369_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT43), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n571_), .A2(new_n629_), .A3(new_n369_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n631_), .A2(KEYINPUT44), .A3(new_n383_), .A4(new_n338_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(new_n573_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n629_), .B1(new_n571_), .B2(new_n369_), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT43), .B(new_n370_), .C1(new_n552_), .C2(new_n570_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n383_), .B(new_n338_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT44), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(G29gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n626_), .B1(new_n633_), .B2(new_n639_), .ZN(G1328gat));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  INV_X1    g440(.A(G36gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n625_), .A2(new_n642_), .A3(new_n589_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT45), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT45), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n625_), .A2(new_n645_), .A3(new_n642_), .A4(new_n589_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n463_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n642_), .B1(new_n648_), .B2(new_n632_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n641_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n646_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n648_), .A2(new_n632_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n651_), .B(KEYINPUT46), .C1(new_n652_), .C2(new_n642_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(G1329gat));
  NAND2_X1  g453(.A1(new_n632_), .A2(new_n604_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n638_), .A2(G43gat), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n579_), .A2(new_n545_), .A3(new_n624_), .ZN(new_n657_));
  OAI22_X1  g456(.A1(new_n655_), .A2(new_n656_), .B1(G43gat), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g458(.A(G50gat), .B1(new_n625_), .B2(new_n620_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n632_), .A2(new_n620_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n638_), .A2(G50gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n661_), .B2(new_n662_), .ZN(G1331gat));
  INV_X1    g462(.A(new_n337_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n571_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n571_), .A2(KEYINPUT103), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n304_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n386_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n669_), .A2(KEYINPUT104), .A3(new_n386_), .A4(new_n670_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n246_), .A4(new_n573_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n670_), .A2(new_n584_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(new_n665_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n573_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G57gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT105), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n675_), .A2(new_n682_), .A3(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1332gat));
  AOI21_X1  g483(.A(new_n247_), .B1(new_n677_), .B2(new_n589_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT48), .Z(new_n686_));
  NOR2_X1   g485(.A1(new_n463_), .A2(G64gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT106), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n673_), .A2(new_n674_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(G1333gat));
  NAND4_X1  g489(.A1(new_n673_), .A2(new_n674_), .A3(new_n253_), .A4(new_n604_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n676_), .A2(new_n665_), .A3(new_n545_), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n692_), .A2(KEYINPUT49), .A3(new_n253_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT49), .B1(new_n692_), .B2(new_n253_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n691_), .A2(KEYINPUT107), .A3(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1334gat));
  AOI21_X1  g499(.A(new_n254_), .B1(new_n677_), .B2(new_n620_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT50), .Z(new_n702_));
  NAND4_X1  g501(.A1(new_n673_), .A2(new_n674_), .A3(new_n254_), .A4(new_n620_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1335gat));
  NAND4_X1  g503(.A1(new_n631_), .A2(new_n383_), .A3(new_n664_), .A4(new_n670_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n705_), .A2(new_n202_), .A3(new_n507_), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n304_), .B(new_n624_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n573_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1336gat));
  NOR3_X1   g508(.A1(new_n705_), .A2(new_n203_), .A3(new_n463_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G92gat), .B1(new_n707_), .B2(new_n589_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1337gat));
  NOR2_X1   g511(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n713_));
  AND2_X1   g512(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n714_));
  OAI21_X1  g513(.A(G99gat), .B1(new_n705_), .B2(new_n545_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n707_), .A2(new_n242_), .A3(new_n604_), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n713_), .B(new_n714_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  AND4_X1   g516(.A1(KEYINPUT108), .A2(new_n715_), .A3(KEYINPUT51), .A4(new_n716_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1338gat));
  XOR2_X1   g518(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n383_), .B(new_n664_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n722_), .A2(new_n304_), .A3(new_n569_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n723_), .B2(new_n219_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n707_), .A2(new_n219_), .A3(new_n620_), .ZN(new_n725_));
  OAI211_X1 g524(.A(G106gat), .B(new_n720_), .C1(new_n705_), .C2(new_n569_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT53), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT53), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n724_), .A2(new_n729_), .A3(new_n726_), .A4(new_n725_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1339gat));
  NAND2_X1  g530(.A1(new_n337_), .A2(new_n297_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT56), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n285_), .A2(new_n282_), .A3(new_n286_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT69), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n281_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT55), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n285_), .A2(new_n282_), .A3(KEYINPUT55), .A4(new_n286_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n281_), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(new_n282_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n285_), .A2(new_n264_), .A3(new_n286_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n276_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n737_), .A2(new_n742_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n733_), .B1(new_n746_), .B2(new_n296_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n740_), .A2(new_n741_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n750_), .A3(new_n744_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n293_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n732_), .B1(new_n747_), .B2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n318_), .A2(new_n319_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n328_), .B2(new_n319_), .ZN(new_n755_));
  MUX2_X1   g554(.A(new_n329_), .B(new_n755_), .S(new_n334_), .Z(new_n756_));
  NAND3_X1  g555(.A1(new_n298_), .A2(new_n299_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT57), .B(new_n582_), .C1(new_n753_), .C2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT112), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n337_), .A2(new_n297_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n293_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n293_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n757_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(KEYINPUT57), .A4(new_n582_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n760_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n582_), .B1(new_n753_), .B2(new_n758_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n756_), .A2(new_n297_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT58), .B(new_n772_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n369_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n771_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n383_), .B1(new_n768_), .B2(new_n778_), .ZN(new_n779_));
  XOR2_X1   g578(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n780_));
  NOR3_X1   g579(.A1(new_n369_), .A2(new_n383_), .A3(new_n337_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n302_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(KEYINPUT110), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n781_), .A2(new_n302_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n782_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n779_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n779_), .A2(KEYINPUT113), .A3(new_n786_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n589_), .A2(new_n507_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n551_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT59), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n760_), .A2(new_n767_), .A3(new_n771_), .A4(new_n777_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n797_), .A2(KEYINPUT114), .A3(new_n383_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT114), .B1(new_n797_), .B2(new_n383_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n785_), .A2(new_n784_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n785_), .B2(new_n780_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n798_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n793_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n796_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n664_), .A2(new_n485_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n779_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n797_), .A2(KEYINPUT114), .A3(new_n383_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n786_), .A3(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n810_), .A2(KEYINPUT115), .A3(new_n803_), .A4(new_n793_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n795_), .A2(new_n805_), .A3(new_n806_), .A4(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n485_), .B1(new_n794_), .B2(new_n664_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(KEYINPUT116), .A3(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1340gat));
  AND3_X1   g617(.A1(new_n789_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n487_), .A2(KEYINPUT60), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n487_), .B1(new_n304_), .B2(KEYINPUT60), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT117), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n795_), .A2(new_n805_), .A3(new_n811_), .ZN(new_n825_));
  OAI21_X1  g624(.A(G120gat), .B1(new_n825_), .B2(new_n304_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1341gat));
  INV_X1    g626(.A(G127gat), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n383_), .A2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n795_), .A2(new_n805_), .A3(new_n811_), .A4(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n794_), .B2(new_n383_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT118), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(new_n834_), .A3(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1342gat));
  XNOR2_X1  g635(.A(KEYINPUT119), .B(G134gat), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n825_), .A2(new_n370_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G134gat), .B1(new_n819_), .B2(new_n583_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1343gat));
  AND2_X1   g639(.A1(new_n789_), .A2(new_n790_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n791_), .A2(new_n550_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT120), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n664_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n469_), .ZN(G1344gat));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n304_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(new_n470_), .ZN(G1345gat));
  NOR2_X1   g647(.A1(new_n844_), .A2(new_n383_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT61), .B(G155gat), .Z(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1346gat));
  NOR3_X1   g650(.A1(new_n844_), .A2(new_n357_), .A3(new_n370_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n841_), .A2(new_n583_), .A3(new_n843_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n357_), .B2(new_n853_), .ZN(G1347gat));
  NOR2_X1   g653(.A1(new_n463_), .A2(new_n573_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n604_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT121), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n620_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n810_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n337_), .A3(new_n397_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n810_), .A2(new_n858_), .A3(new_n337_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n863_), .A2(G169gat), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n864_), .A2(new_n865_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n862_), .A2(new_n866_), .A3(new_n867_), .ZN(G1348gat));
  NAND2_X1  g667(.A1(new_n861_), .A2(new_n670_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n841_), .A2(new_n858_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n304_), .A2(new_n398_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n869_), .A2(new_n398_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  AOI21_X1  g671(.A(G183gat), .B1(new_n870_), .B2(new_n384_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n859_), .B(KEYINPUT123), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n383_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n407_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n875_), .B2(new_n876_), .ZN(G1350gat));
  OAI21_X1  g676(.A(G190gat), .B1(new_n874_), .B2(new_n370_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n861_), .A2(new_n583_), .A3(new_n408_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1351gat));
  NAND4_X1  g679(.A1(new_n789_), .A2(new_n550_), .A3(new_n790_), .A4(new_n855_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n664_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(new_n333_), .ZN(G1352gat));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n304_), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(G204gat), .Z(G1353gat));
  AOI21_X1  g684(.A(new_n383_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT124), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n881_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n889_));
  OR3_X1    g688(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n888_), .B2(new_n890_), .ZN(G1354gat));
  XNOR2_X1  g691(.A(KEYINPUT127), .B(G218gat), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n881_), .A2(new_n370_), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895_));
  OR3_X1    g694(.A1(new_n881_), .A2(new_n895_), .A3(new_n582_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n881_), .B2(new_n582_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n894_), .B1(new_n898_), .B2(new_n893_), .ZN(G1355gat));
endmodule


