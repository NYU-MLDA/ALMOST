//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  AND2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT85), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n207_), .B1(new_n211_), .B2(KEYINPUT86), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n210_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT86), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  AOI211_X1 g014(.A(new_n204_), .B(new_n205_), .C1(new_n212_), .C2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n204_), .A2(KEYINPUT2), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n205_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n204_), .A2(KEYINPUT2), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n222_), .A2(new_n209_), .A3(new_n206_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n216_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT84), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n226_), .B(new_n227_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n228_), .B1(new_n229_), .B2(new_n225_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT99), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n216_), .A2(new_n223_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n231_), .A2(KEYINPUT98), .B1(new_n236_), .B2(new_n229_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT98), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n224_), .A2(new_n238_), .A3(new_n230_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n237_), .A2(new_n239_), .B1(KEYINPUT99), .B2(new_n232_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n203_), .B(new_n235_), .C1(new_n240_), .C2(new_n234_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G1gat), .B(G29gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G85gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G57gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n202_), .A3(new_n239_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT100), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n241_), .A2(KEYINPUT100), .A3(new_n245_), .A4(new_n246_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n246_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n245_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n250_), .A3(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G197gat), .B(G204gat), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT89), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(KEYINPUT21), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(KEYINPUT21), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT88), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n257_), .B1(new_n255_), .B2(KEYINPUT21), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT91), .Z(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT23), .ZN(new_n266_));
  INV_X1    g065(.A(G169gat), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n266_), .B1(KEYINPUT24), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT93), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n269_), .A2(KEYINPUT24), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT25), .B(G183gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n271_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT22), .B(G169gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n268_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n272_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n266_), .B1(G183gat), .B2(G190gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n264_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT20), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(KEYINPUT82), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n281_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n283_), .A3(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n270_), .A2(new_n273_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n277_), .B(KEYINPUT81), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n287_), .B1(new_n294_), .B2(new_n263_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n286_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n284_), .B(KEYINPUT94), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n278_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n263_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT20), .B1(new_n294_), .B2(new_n263_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n299_), .B1(new_n300_), .B2(KEYINPUT92), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(KEYINPUT92), .B2(new_n300_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G226gat), .A2(G233gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT19), .Z(new_n304_));
  MUX2_X1   g103(.A(new_n296_), .B(new_n302_), .S(new_n304_), .Z(new_n305_));
  XOR2_X1   g104(.A(G64gat), .B(G92gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT97), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT96), .B(KEYINPUT18), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G8gat), .B(G36gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n305_), .A2(KEYINPUT32), .A3(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n295_), .B(new_n304_), .C1(new_n263_), .C2(new_n298_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n315_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n302_), .A2(new_n304_), .ZN(new_n319_));
  AOI211_X1 g118(.A(new_n318_), .B(new_n319_), .C1(KEYINPUT32), .C2(new_n312_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n313_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n247_), .A2(KEYINPUT33), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT33), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n241_), .A2(new_n323_), .A3(new_n245_), .A4(new_n246_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n237_), .A2(new_n203_), .A3(new_n239_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n252_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n235_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n240_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(KEYINPUT4), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(new_n330_), .B2(new_n202_), .ZN(new_n331_));
  OR3_X1    g130(.A1(new_n319_), .A2(new_n318_), .A3(new_n311_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n311_), .B1(new_n319_), .B2(new_n318_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n254_), .A2(new_n321_), .B1(new_n325_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(G228gat), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n340_), .B(new_n263_), .C1(new_n236_), .C2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n345_));
  NAND2_X1  g144(.A1(new_n224_), .A2(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n346_), .A2(new_n264_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n342_), .B(new_n344_), .C1(new_n347_), .C2(new_n340_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n340_), .B1(new_n346_), .B2(new_n264_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n342_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n343_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n236_), .A2(new_n341_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n353_), .B(KEYINPUT28), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n352_), .A2(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n348_), .A2(new_n358_), .A3(new_n360_), .A4(new_n351_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT83), .B(G43gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n294_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(new_n230_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(G15gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT30), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT31), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n369_), .B(new_n374_), .Z(new_n375_));
  NAND2_X1  g174(.A1(new_n364_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n364_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n362_), .A2(new_n375_), .A3(new_n363_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n305_), .A2(new_n311_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n332_), .A3(KEYINPUT27), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT101), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n334_), .B2(new_n384_), .ZN(new_n385_));
  AOI211_X1 g184(.A(KEYINPUT101), .B(KEYINPUT27), .C1(new_n332_), .C2(new_n333_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n380_), .B(new_n382_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  OAI22_X1  g186(.A1(new_n336_), .A2(new_n376_), .B1(new_n387_), .B2(new_n254_), .ZN(new_n388_));
  INV_X1    g187(.A(G85gat), .ZN(new_n389_));
  INV_X1    g188(.A(G92gat), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n389_), .A2(new_n390_), .A3(KEYINPUT9), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n392_));
  AND3_X1   g191(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G85gat), .B(G92gat), .Z(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT9), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT64), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT10), .B(G99gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G106gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n398_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n394_), .B(new_n396_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT8), .ZN(new_n404_));
  INV_X1    g203(.A(G99gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n400_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT7), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(KEYINPUT65), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT65), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(KEYINPUT7), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n406_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT66), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n393_), .B2(new_n392_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G99gat), .A2(G106gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(KEYINPUT66), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n409_), .A2(KEYINPUT7), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n405_), .A3(new_n400_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n411_), .A2(new_n413_), .A3(new_n418_), .A4(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n404_), .B1(new_n421_), .B2(new_n395_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n395_), .A2(new_n404_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n407_), .A2(KEYINPUT65), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n419_), .A2(new_n424_), .B1(new_n405_), .B2(new_n400_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n408_), .A2(new_n406_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n393_), .A2(new_n392_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n423_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n403_), .B1(new_n422_), .B2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G29gat), .B(G36gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G43gat), .B(G50gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT15), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G232gat), .A2(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT34), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n437_), .A2(KEYINPUT35), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n438_), .A2(KEYINPUT73), .ZN(new_n439_));
  INV_X1    g238(.A(new_n433_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n435_), .B(new_n439_), .C1(new_n440_), .C2(new_n430_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(KEYINPUT35), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G190gat), .B(G218gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(G134gat), .B(G162gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT36), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n443_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n443_), .A2(KEYINPUT72), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n449_), .A2(KEYINPUT36), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n443_), .A2(KEYINPUT72), .A3(new_n453_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n451_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n388_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G230gat), .A2(G233gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n462_), .A2(new_n463_), .A3(G78gat), .ZN(new_n464_));
  INV_X1    g263(.A(G78gat), .ZN(new_n465_));
  OR2_X1    g264(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(new_n461_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n460_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G57gat), .B(G64gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(G78gat), .B1(new_n462_), .B2(new_n463_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n465_), .A3(new_n461_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT11), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n469_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n474_), .A2(new_n470_), .A3(KEYINPUT11), .A4(new_n471_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n430_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n475_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n478_), .B(new_n403_), .C1(new_n422_), .C2(new_n429_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n459_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n477_), .A2(new_n479_), .B1(new_n481_), .B2(new_n430_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n477_), .B2(new_n485_), .ZN(new_n486_));
  AOI211_X1 g285(.A(KEYINPUT69), .B(new_n484_), .C1(new_n430_), .C2(new_n476_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n482_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n480_), .B1(new_n488_), .B2(new_n459_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G120gat), .B(G148gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT5), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n489_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n496_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G1gat), .B(G8gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT74), .ZN(new_n501_));
  INV_X1    g300(.A(G22gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n371_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G15gat), .A2(G22gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G1gat), .A2(G8gat), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n503_), .A2(new_n504_), .B1(KEYINPUT14), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n501_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n434_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n500_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(new_n506_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n433_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n508_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT78), .ZN(new_n515_));
  INV_X1    g314(.A(new_n513_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n507_), .A2(new_n440_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n511_), .A2(new_n433_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT77), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n507_), .A2(new_n440_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n512_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(KEYINPUT77), .A3(new_n516_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  AND3_X1   g327(.A1(new_n515_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n515_), .B2(new_n525_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT79), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n515_), .A2(new_n525_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n515_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT79), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n532_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n499_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n478_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(new_n507_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G127gat), .B(G155gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT16), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G183gat), .B(G211gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  MUX2_X1   g348(.A(new_n545_), .B(KEYINPUT17), .S(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(KEYINPUT75), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT76), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n550_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n540_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n458_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n254_), .ZN(new_n558_));
  OAI21_X1  g357(.A(G1gat), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT103), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT103), .B(G1gat), .C1(new_n557_), .C2(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT80), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n538_), .A2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT80), .B1(new_n532_), .B2(new_n537_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n388_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n457_), .A2(new_n570_), .ZN(new_n571_));
  AOI211_X1 g370(.A(KEYINPUT37), .B(new_n451_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n574_), .A2(new_n555_), .A3(new_n499_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n569_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT102), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT102), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n569_), .A2(new_n578_), .A3(new_n575_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n558_), .A2(G1gat), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n577_), .A2(KEYINPUT38), .A3(new_n579_), .A4(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT38), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n563_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT104), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n563_), .A2(new_n584_), .A3(KEYINPUT104), .A4(new_n581_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(G1324gat));
  OR2_X1    g388(.A1(new_n385_), .A2(new_n386_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n382_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G8gat), .B1(new_n557_), .B2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT39), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT39), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n577_), .A2(new_n579_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n592_), .A2(G8gat), .ZN(new_n597_));
  OAI22_X1  g396(.A1(new_n594_), .A2(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  OAI221_X1 g400(.A(new_n599_), .B1(new_n596_), .B2(new_n597_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1325gat));
  INV_X1    g402(.A(new_n596_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G15gat), .B1(new_n557_), .B2(new_n375_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n608_), .A3(new_n609_), .ZN(G1326gat));
  OAI21_X1  g409(.A(G22gat), .B1(new_n557_), .B2(new_n364_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT42), .ZN(new_n612_));
  INV_X1    g411(.A(new_n364_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n604_), .A2(new_n502_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(G1327gat));
  NOR3_X1   g414(.A1(new_n499_), .A2(new_n554_), .A3(new_n457_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n569_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(G29gat), .B1(new_n618_), .B2(new_n254_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n540_), .A2(new_n554_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT43), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n388_), .A2(new_n621_), .A3(new_n574_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n388_), .B2(new_n574_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n620_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT44), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n626_), .A2(G29gat), .A3(new_n254_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n623_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n388_), .A2(new_n621_), .A3(new_n574_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(KEYINPUT44), .A3(new_n620_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n619_), .B1(new_n627_), .B2(new_n631_), .ZN(G1328gat));
  INV_X1    g431(.A(G36gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n592_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n634_), .B2(new_n631_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n569_), .A2(new_n633_), .A3(new_n591_), .A4(new_n616_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT45), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(KEYINPUT46), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT46), .ZN(new_n640_));
  INV_X1    g439(.A(new_n638_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(new_n635_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(G1329gat));
  NAND3_X1  g442(.A1(new_n569_), .A2(new_n377_), .A3(new_n616_), .ZN(new_n644_));
  INV_X1    g443(.A(G43gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(KEYINPUT107), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n626_), .A2(G43gat), .A3(new_n377_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n631_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT47), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT47), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n650_), .B(new_n655_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1330gat));
  OR3_X1    g456(.A1(new_n617_), .A2(G50gat), .A3(new_n364_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n631_), .A2(new_n626_), .A3(new_n613_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT108), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n659_), .A2(new_n660_), .A3(G50gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n659_), .B2(G50gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(G1331gat));
  INV_X1    g462(.A(new_n499_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n568_), .A2(new_n664_), .A3(new_n555_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n458_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G57gat), .B1(new_n667_), .B2(new_n558_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n388_), .A2(new_n538_), .ZN(new_n669_));
  AND4_X1   g468(.A1(new_n499_), .A2(new_n669_), .A3(new_n554_), .A4(new_n573_), .ZN(new_n670_));
  INV_X1    g469(.A(G57gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n671_), .A3(new_n254_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n668_), .A2(new_n672_), .ZN(G1332gat));
  INV_X1    g472(.A(G64gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n666_), .B2(new_n591_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT48), .Z(new_n676_));
  NAND3_X1  g475(.A1(new_n670_), .A2(new_n674_), .A3(new_n591_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1333gat));
  INV_X1    g477(.A(G71gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n666_), .B2(new_n377_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT49), .Z(new_n681_));
  NAND3_X1  g480(.A1(new_n670_), .A2(new_n679_), .A3(new_n377_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1334gat));
  AOI21_X1  g482(.A(new_n465_), .B1(new_n666_), .B2(new_n613_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT50), .Z(new_n685_));
  NAND3_X1  g484(.A1(new_n670_), .A2(new_n465_), .A3(new_n613_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1335gat));
  INV_X1    g486(.A(new_n538_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n664_), .A2(new_n554_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n630_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G85gat), .B1(new_n690_), .B2(new_n558_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n457_), .ZN(new_n692_));
  AND4_X1   g491(.A1(new_n499_), .A2(new_n669_), .A3(new_n555_), .A4(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n389_), .A3(new_n254_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1336gat));
  OAI21_X1  g494(.A(G92gat), .B1(new_n690_), .B2(new_n592_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n390_), .A3(new_n591_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1337gat));
  OAI21_X1  g497(.A(G99gat), .B1(new_n690_), .B2(new_n375_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n693_), .A2(new_n377_), .A3(new_n399_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g501(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n613_), .B(new_n689_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G106gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT52), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n707_), .A3(G106gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n693_), .A2(new_n400_), .A3(new_n613_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n703_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n704_), .A2(new_n707_), .A3(G106gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n704_), .B2(G106gat), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n710_), .B(new_n703_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n711_), .A2(new_n715_), .ZN(G1339gat));
  NAND2_X1  g515(.A1(new_n489_), .A2(new_n494_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n531_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n535_), .A2(KEYINPUT79), .A3(new_n536_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n477_), .A2(new_n479_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n430_), .A2(new_n481_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n477_), .A2(new_n485_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT69), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n477_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n724_), .A2(new_n726_), .A3(new_n459_), .A4(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT110), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT55), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(KEYINPUT110), .A3(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT111), .B1(new_n488_), .B2(new_n459_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(G230gat), .A4(G233gat), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n730_), .A2(new_n732_), .A3(new_n733_), .A4(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n493_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT56), .B1(new_n737_), .B2(new_n493_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n721_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n523_), .A2(new_n513_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n508_), .A2(new_n512_), .A3(new_n516_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n534_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n742_), .B1(new_n536_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n536_), .A2(new_n742_), .A3(new_n745_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n495_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n692_), .B1(new_n741_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT57), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT57), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n717_), .B1(new_n532_), .B2(new_n537_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n737_), .A2(new_n493_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n754_), .B1(new_n757_), .B2(new_n738_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n750_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n457_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n748_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n717_), .B1(new_n761_), .B2(new_n746_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n757_), .B2(new_n738_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n573_), .B1(new_n763_), .B2(KEYINPUT58), .ZN(new_n764_));
  INV_X1    g563(.A(new_n762_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT113), .B(KEYINPUT58), .Z(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n753_), .A2(new_n760_), .B1(new_n764_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n752_), .B1(new_n770_), .B2(KEYINPUT115), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n765_), .B(KEYINPUT58), .C1(new_n739_), .C2(new_n740_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n574_), .C1(new_n763_), .C2(new_n767_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(KEYINPUT115), .C1(KEYINPUT57), .C2(new_n751_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n555_), .B1(new_n771_), .B2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n664_), .A2(new_n554_), .A3(new_n567_), .A4(new_n573_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT54), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n591_), .A2(new_n558_), .A3(new_n378_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n554_), .B1(new_n770_), .B2(new_n752_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n777_), .B(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n784_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n773_), .B1(KEYINPUT57), .B2(new_n751_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n752_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n555_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT114), .A3(new_n778_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n788_), .A2(new_n792_), .A3(new_n780_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n783_), .B1(new_n793_), .B2(new_n781_), .ZN(new_n794_));
  OAI21_X1  g593(.A(G113gat), .B1(new_n794_), .B2(new_n567_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n788_), .A2(new_n792_), .A3(new_n780_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n797_), .A2(G113gat), .A3(new_n538_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(new_n796_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(G113gat), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n797_), .A2(KEYINPUT59), .B1(new_n779_), .B2(new_n782_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n568_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT116), .B1(new_n803_), .B2(new_n798_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n804_), .ZN(G1340gat));
  OAI21_X1  g604(.A(G120gat), .B1(new_n794_), .B2(new_n664_), .ZN(new_n806_));
  INV_X1    g605(.A(G120gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n664_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(KEYINPUT60), .B2(new_n807_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n806_), .B1(new_n797_), .B2(new_n809_), .ZN(G1341gat));
  AOI21_X1  g609(.A(G127gat), .B1(new_n793_), .B2(new_n554_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n554_), .A2(G127gat), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(KEYINPUT117), .Z(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n802_), .B2(new_n813_), .ZN(G1342gat));
  AOI21_X1  g613(.A(G134gat), .B1(new_n793_), .B2(new_n692_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n574_), .A2(G134gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT118), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n802_), .B2(new_n817_), .ZN(G1343gat));
  NAND2_X1  g617(.A1(new_n788_), .A2(new_n792_), .ZN(new_n819_));
  NOR4_X1   g618(.A1(new_n819_), .A2(new_n558_), .A3(new_n379_), .A4(new_n591_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n688_), .ZN(new_n821_));
  XOR2_X1   g620(.A(KEYINPUT119), .B(G141gat), .Z(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1344gat));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n499_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n554_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1346gat));
  AOI21_X1  g627(.A(G162gat), .B1(new_n820_), .B2(new_n692_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n574_), .A2(G162gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT120), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n820_), .B2(new_n831_), .ZN(G1347gat));
  NOR3_X1   g631(.A1(new_n592_), .A2(new_n254_), .A3(new_n375_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n364_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n267_), .B1(new_n835_), .B2(new_n688_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n836_), .A2(KEYINPUT62), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(KEYINPUT62), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n279_), .A3(new_n688_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(G1348gat));
  NAND3_X1  g639(.A1(new_n833_), .A2(G176gat), .A3(new_n499_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n788_), .A2(new_n364_), .A3(new_n792_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n788_), .A2(new_n792_), .A3(KEYINPUT121), .A4(new_n364_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847_));
  AOI21_X1  g646(.A(G176gat), .B1(new_n835_), .B2(new_n499_), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1349gat));
  NOR2_X1   g650(.A1(new_n555_), .A2(new_n275_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n835_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n833_), .A2(new_n554_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n855_), .B2(G183gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT123), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n853_), .B(new_n858_), .C1(new_n855_), .C2(G183gat), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1350gat));
  NAND2_X1  g659(.A1(new_n835_), .A2(new_n574_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G190gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n835_), .A2(new_n276_), .A3(new_n692_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1351gat));
  AND2_X1   g663(.A1(new_n788_), .A2(new_n792_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n592_), .A2(new_n254_), .A3(new_n379_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n867_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n688_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n865_), .A2(new_n688_), .A3(new_n866_), .ZN(new_n870_));
  INV_X1    g669(.A(G197gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n871_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n868_), .A2(new_n872_), .A3(new_n873_), .ZN(G1352gat));
  NAND2_X1  g673(.A1(new_n867_), .A2(new_n499_), .ZN(new_n875_));
  OR2_X1    g674(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT126), .Z(new_n878_));
  AND3_X1   g677(.A1(new_n875_), .A2(new_n876_), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1353gat));
  XOR2_X1   g680(.A(KEYINPUT63), .B(G211gat), .Z(new_n882_));
  AND3_X1   g681(.A1(new_n867_), .A2(new_n554_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n867_), .A2(new_n554_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1354gat));
  AOI21_X1  g685(.A(G218gat), .B1(new_n867_), .B2(new_n692_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n574_), .A2(G218gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT127), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n867_), .B2(new_n889_), .ZN(G1355gat));
endmodule


