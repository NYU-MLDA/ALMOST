//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n202_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(KEYINPUT21), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT82), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT82), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G155gat), .A3(G162gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n209_), .B1(new_n214_), .B2(KEYINPUT1), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n211_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT83), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT83), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n211_), .A2(new_n213_), .A3(new_n219_), .A4(new_n216_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n215_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G141gat), .B(G148gat), .Z(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n209_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n212_), .B1(G155gat), .B2(G162gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n210_), .A2(KEYINPUT82), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n214_), .A2(KEYINPUT86), .A3(new_n224_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT85), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G141gat), .A2(G148gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n236_), .A2(KEYINPUT84), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT84), .B1(new_n236_), .B2(new_n237_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n235_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n229_), .B(new_n230_), .C1(new_n232_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n223_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n244_));
  OAI21_X1  g043(.A(new_n208_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G228gat), .A3(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G78gat), .B(G106gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n242_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n223_), .A2(new_n241_), .A3(KEYINPUT87), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT29), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G228gat), .A2(G233gat), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n208_), .A2(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n252_), .A2(KEYINPUT88), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT88), .B1(new_n252_), .B2(new_n254_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n246_), .B(new_n248_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT90), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n246_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n247_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n223_), .A2(new_n241_), .A3(KEYINPUT87), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT87), .B1(new_n223_), .B2(new_n241_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT29), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n254_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n262_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n252_), .A2(KEYINPUT88), .A3(new_n254_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n270_), .A2(KEYINPUT90), .A3(new_n246_), .A4(new_n248_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT29), .B1(new_n250_), .B2(new_n251_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G22gat), .B(G50gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT28), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n272_), .A2(new_n274_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n259_), .A2(new_n261_), .A3(new_n271_), .A4(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT91), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n260_), .B2(new_n247_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT91), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n282_), .A2(new_n259_), .A3(new_n283_), .A4(new_n271_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G15gat), .B(G43gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n288_), .A2(KEYINPUT24), .ZN(new_n289_));
  INV_X1    g088(.A(G183gat), .ZN(new_n290_));
  INV_X1    g089(.A(G190gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT23), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n288_), .A2(KEYINPUT24), .A3(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n289_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n290_), .A2(KEYINPUT76), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G183gat), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n300_), .A2(new_n302_), .A3(KEYINPUT25), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G183gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n303_), .A2(new_n309_), .A3(KEYINPUT77), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311_));
  INV_X1    g110(.A(new_n308_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n312_), .A2(new_n306_), .B1(new_n304_), .B2(G183gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n300_), .A2(new_n302_), .A3(KEYINPUT25), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n299_), .B1(new_n310_), .B2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n300_), .A2(new_n302_), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n317_), .A2(new_n291_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT22), .B(G169gat), .ZN(new_n319_));
  INV_X1    g118(.A(G176gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n296_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT78), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT77), .B1(new_n303_), .B2(new_n309_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n313_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n298_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n318_), .A2(new_n322_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT78), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n330_), .A3(KEYINPUT30), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT30), .B1(new_n325_), .B2(new_n330_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G227gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n332_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n325_), .A2(new_n330_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT30), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n338_), .B1(new_n341_), .B2(new_n331_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n287_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n336_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n331_), .A3(new_n338_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n286_), .A3(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n344_), .A3(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G113gat), .B(G120gat), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n350_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT79), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n348_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n348_), .A2(new_n359_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n344_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n261_), .A2(new_n257_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n278_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n285_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT0), .ZN(new_n369_));
  INV_X1    g168(.A(G57gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G85gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n250_), .A2(new_n251_), .A3(new_n356_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n351_), .A2(new_n353_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n243_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(KEYINPUT4), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT97), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n374_), .A2(KEYINPUT97), .A3(KEYINPUT4), .A4(new_n376_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n374_), .A2(KEYINPUT4), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n374_), .A2(new_n376_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n387_), .A2(new_n385_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n373_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n381_), .B1(new_n378_), .B2(new_n377_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n384_), .A3(new_n380_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n372_), .B1(new_n387_), .B2(new_n385_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT33), .B1(new_n390_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n339_), .A2(new_n208_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n295_), .B1(G183gat), .B2(G190gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n296_), .B(KEYINPUT95), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n399_), .A2(new_n321_), .A3(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n402_));
  INV_X1    g201(.A(new_n288_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n402_), .A2(new_n403_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(new_n288_), .A3(new_n296_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT92), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n312_), .A2(new_n408_), .A3(new_n306_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT92), .B1(new_n307_), .B2(new_n308_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT25), .B(G183gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT94), .B1(new_n407_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT94), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n404_), .A2(new_n412_), .A3(new_n415_), .A4(new_n406_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n401_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n206_), .B(new_n207_), .Z(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT20), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n397_), .B1(new_n398_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n397_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT20), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n339_), .A2(new_n208_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT96), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n420_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G8gat), .B(G36gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT18), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G64gat), .ZN(new_n431_));
  INV_X1    g230(.A(G92gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n428_), .A2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n420_), .B(new_n433_), .C1(new_n426_), .C2(new_n427_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n384_), .B1(new_n391_), .B2(new_n380_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n372_), .B1(new_n438_), .B2(new_n388_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n433_), .A2(KEYINPUT32), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n428_), .A2(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n398_), .A2(new_n419_), .A3(new_n397_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT98), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n208_), .A2(new_n401_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n407_), .A2(new_n413_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT20), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n418_), .B1(new_n325_), .B2(new_n330_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n397_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n444_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n450_), .A2(new_n445_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n443_), .B1(new_n453_), .B2(new_n442_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n386_), .A2(new_n373_), .A3(new_n389_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n439_), .A2(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n395_), .A2(new_n441_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n367_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n285_), .A2(new_n366_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n364_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n362_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n363_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n360_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n285_), .A2(new_n463_), .A3(new_n366_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n466_), .B1(new_n453_), .B2(new_n434_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT99), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n436_), .A2(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n436_), .A2(new_n468_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n437_), .A2(new_n466_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n456_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n458_), .B1(new_n465_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G190gat), .B(G218gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G134gat), .B(G162gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n478_), .B(KEYINPUT36), .Z(new_n479_));
  NAND2_X1  g278(.A1(G232gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT34), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(KEYINPUT35), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT10), .B(G99gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT64), .ZN(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G85gat), .B(G92gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT65), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT9), .ZN(new_n490_));
  INV_X1    g289(.A(G85gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(new_n432_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n487_), .A2(new_n488_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT8), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT7), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n486_), .A2(new_n493_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT6), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n487_), .A2(KEYINPUT8), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n496_), .A2(new_n499_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n487_), .A2(KEYINPUT8), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G29gat), .B(G36gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT15), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n482_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n481_), .A2(KEYINPUT35), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n512_), .B(KEYINPUT69), .Z(new_n513_));
  NAND3_X1  g312(.A1(new_n501_), .A2(new_n509_), .A3(new_n505_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n514_), .A2(new_n515_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n511_), .B(new_n513_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n514_), .B(new_n515_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n513_), .B1(new_n520_), .B2(new_n511_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n479_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT71), .ZN(new_n523_));
  INV_X1    g322(.A(new_n521_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n478_), .A2(KEYINPUT36), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n518_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT71), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n527_), .B(new_n479_), .C1(new_n519_), .C2(new_n521_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n523_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT37), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n526_), .A2(new_n522_), .A3(KEYINPUT37), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n475_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G71gat), .B(G78gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(KEYINPUT11), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  AND3_X1   g338(.A1(new_n501_), .A2(new_n505_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n539_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n541_));
  OAI22_X1  g340(.A1(new_n540_), .A2(new_n541_), .B1(KEYINPUT66), .B2(KEYINPUT12), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT66), .B(KEYINPUT12), .Z(new_n543_));
  OR2_X1    g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G230gat), .A2(G233gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(G230gat), .B(G233gat), .C1(new_n540_), .C2(new_n541_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G120gat), .B(G148gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G204gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT5), .B(G176gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n552_), .B(KEYINPUT67), .Z(new_n555_));
  OAI211_X1 g354(.A(new_n553_), .B(new_n554_), .C1(new_n548_), .C2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n553_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n548_), .A2(new_n555_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n560_));
  OAI21_X1  g359(.A(new_n556_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G15gat), .B(G22gat), .Z(new_n562_));
  NAND2_X1  g361(.A1(G1gat), .A2(G8gat), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(KEYINPUT14), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT72), .ZN(new_n565_));
  XOR2_X1   g364(.A(G1gat), .B(G8gat), .Z(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(new_n509_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n567_), .A2(new_n568_), .A3(new_n510_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n569_), .B2(new_n509_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n570_), .A2(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(G197gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT75), .B(G169gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n575_), .A2(new_n579_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n561_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G183gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(G211gat), .Z(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT17), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT73), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(KEYINPUT17), .B2(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n569_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n539_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n590_), .A2(KEYINPUT74), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(KEYINPUT73), .B2(new_n589_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n593_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n597_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n584_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n534_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n534_), .A2(KEYINPUT100), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT101), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n607_), .A2(new_n611_), .A3(new_n608_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n456_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(G1gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT38), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n610_), .A2(KEYINPUT38), .A3(new_n612_), .A4(new_n614_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n529_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n475_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n604_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n613_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1324gat));
  NAND2_X1  g424(.A1(new_n610_), .A2(new_n612_), .ZN(new_n626_));
  INV_X1    g425(.A(G8gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n473_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n620_), .A2(new_n604_), .A3(new_n473_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n629_), .A2(KEYINPUT103), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n627_), .B1(new_n629_), .B2(KEYINPUT103), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n634_));
  OAI22_X1  g433(.A1(new_n626_), .A2(new_n628_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT40), .Z(G1325gat));
  NOR3_X1   g435(.A1(new_n609_), .A2(G15gat), .A3(new_n364_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT105), .Z(new_n638_));
  OAI21_X1  g437(.A(G15gat), .B1(new_n621_), .B2(new_n364_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT41), .Z(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n638_), .A2(new_n642_), .A3(new_n643_), .ZN(G1326gat));
  INV_X1    g443(.A(new_n459_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G22gat), .B1(new_n621_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT42), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n645_), .A2(G22gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n609_), .B2(new_n648_), .ZN(G1327gat));
  INV_X1    g448(.A(G29gat), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  INV_X1    g450(.A(new_n532_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n285_), .A2(new_n463_), .A3(new_n366_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n463_), .B1(new_n285_), .B2(new_n366_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n474_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n367_), .A2(new_n457_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n651_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT106), .B(KEYINPUT43), .C1(new_n475_), .C2(new_n653_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n659_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n584_), .A2(new_n602_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(KEYINPUT44), .A3(new_n664_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n456_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n650_), .B1(new_n670_), .B2(KEYINPUT107), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n671_), .B1(KEYINPUT107), .B2(new_n670_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n475_), .A2(new_n529_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n664_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n650_), .A3(new_n456_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n672_), .A2(new_n676_), .ZN(G1328gat));
  NAND2_X1  g476(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n673_), .A2(new_n680_), .A3(new_n473_), .A4(new_n664_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(KEYINPUT45), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(KEYINPUT45), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n667_), .A2(new_n473_), .A3(new_n668_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n680_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n667_), .A2(KEYINPUT108), .A3(new_n473_), .A4(new_n668_), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n679_), .B(new_n686_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n687_), .A2(new_n688_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(G36gat), .A3(new_n690_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n686_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n678_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n691_), .A2(new_n695_), .ZN(G1329gat));
  INV_X1    g495(.A(G43gat), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n364_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n667_), .A2(new_n668_), .A3(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n674_), .B2(new_n364_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT110), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n699_), .A2(new_n703_), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n702_), .A2(KEYINPUT47), .A3(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n675_), .B2(new_n459_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n459_), .A2(G50gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n669_), .B2(new_n711_), .ZN(G1331gat));
  INV_X1    g511(.A(new_n561_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n582_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n603_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n620_), .A2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT111), .Z(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n613_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n534_), .A2(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n456_), .A2(new_n370_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(G1332gat));
  INV_X1    g520(.A(new_n473_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G64gat), .B1(new_n717_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n722_), .A2(G64gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n719_), .B2(new_n726_), .ZN(G1333gat));
  OR3_X1    g526(.A1(new_n719_), .A2(G71gat), .A3(new_n364_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G71gat), .B1(new_n717_), .B2(new_n364_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n729_), .A2(new_n730_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n717_), .B2(new_n645_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n645_), .A2(G78gat), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT114), .Z(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n719_), .B2(new_n737_), .ZN(G1335gat));
  NOR2_X1   g537(.A1(new_n714_), .A2(new_n602_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n663_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n613_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n673_), .A2(new_n739_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n491_), .A3(new_n456_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1336gat));
  OAI21_X1  g543(.A(G92gat), .B1(new_n740_), .B2(new_n722_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n432_), .A3(new_n473_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1337gat));
  INV_X1    g546(.A(KEYINPUT115), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n663_), .A2(new_n463_), .A3(new_n739_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n463_), .A2(new_n484_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n749_), .A2(G99gat), .B1(new_n742_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT51), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n751_), .B2(new_n748_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n753_), .B2(new_n756_), .ZN(G1338gat));
  AOI21_X1  g556(.A(new_n485_), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n740_), .B2(new_n645_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n742_), .A2(new_n485_), .A3(new_n459_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n760_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g564(.A(KEYINPUT121), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n545_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n546_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n542_), .A2(new_n544_), .A3(KEYINPUT55), .A4(new_n545_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n555_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n553_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n569_), .A2(new_n509_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n774_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n579_), .B(new_n775_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n580_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT56), .B(new_n555_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n773_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n533_), .B1(new_n780_), .B2(KEYINPUT58), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n769_), .A2(new_n770_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n555_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n771_), .A2(new_n772_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n785_), .A2(new_n553_), .A3(new_n777_), .A4(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT120), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n780_), .A2(new_n790_), .A3(KEYINPUT58), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n781_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n773_), .A2(new_n582_), .A3(new_n779_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n777_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n529_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n785_), .A2(new_n583_), .A3(new_n553_), .A4(new_n786_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n619_), .B1(new_n799_), .B2(new_n794_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(KEYINPUT57), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n792_), .A2(new_n798_), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n766_), .B1(new_n802_), .B2(new_n602_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n603_), .A2(new_n583_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n653_), .A2(new_n805_), .A3(new_n561_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT118), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(KEYINPUT118), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n804_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n806_), .A2(KEYINPUT118), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT54), .A3(new_n807_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n789_), .A2(new_n791_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n653_), .B1(new_n788_), .B2(new_n787_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n815_), .A2(new_n816_), .B1(KEYINPUT57), .B2(new_n800_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n801_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(KEYINPUT121), .A3(new_n603_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n803_), .A2(new_n814_), .A3(new_n820_), .ZN(new_n821_));
  NOR4_X1   g620(.A1(new_n464_), .A2(new_n473_), .A3(KEYINPUT59), .A4(new_n613_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n464_), .A2(new_n613_), .A3(new_n473_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n800_), .B2(KEYINPUT57), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n796_), .A2(KEYINPUT119), .A3(new_n797_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n602_), .B1(new_n827_), .B2(new_n817_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n823_), .B1(new_n828_), .B2(new_n813_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n821_), .A2(new_n822_), .B1(new_n829_), .B2(KEYINPUT59), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n583_), .A2(G113gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(KEYINPUT122), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(KEYINPUT122), .ZN(new_n833_));
  INV_X1    g632(.A(new_n829_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n583_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1340gat));
  INV_X1    g635(.A(new_n830_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G120gat), .B1(new_n837_), .B2(new_n561_), .ZN(new_n838_));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT60), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n561_), .B2(KEYINPUT60), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(KEYINPUT123), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(KEYINPUT123), .B2(new_n841_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n829_), .B2(new_n843_), .ZN(G1341gat));
  INV_X1    g643(.A(G127gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n830_), .B2(new_n602_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n829_), .A2(G127gat), .A3(new_n603_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT124), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n821_), .A2(new_n822_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n602_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G127gat), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853_));
  INV_X1    g652(.A(new_n847_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n848_), .A2(new_n855_), .ZN(G1342gat));
  OAI21_X1  g655(.A(G134gat), .B1(new_n837_), .B2(new_n653_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n529_), .A2(G134gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n829_), .B2(new_n858_), .ZN(G1343gat));
  NOR2_X1   g658(.A1(new_n828_), .A2(new_n813_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n460_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n456_), .A3(new_n722_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n582_), .ZN(new_n863_));
  INV_X1    g662(.A(G141gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1344gat));
  NOR2_X1   g664(.A1(new_n862_), .A2(new_n561_), .ZN(new_n866_));
  INV_X1    g665(.A(G148gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1345gat));
  NOR2_X1   g667(.A1(new_n862_), .A2(new_n603_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT61), .B(G155gat), .Z(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n862_), .B2(new_n653_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n529_), .A2(G162gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n862_), .B2(new_n873_), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n722_), .A2(new_n456_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n463_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n459_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n821_), .A2(new_n583_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G169gat), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n821_), .A2(new_n877_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n583_), .A3(new_n319_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n881_), .A2(new_n882_), .A3(new_n884_), .ZN(G1348gat));
  OAI21_X1  g684(.A(new_n645_), .B1(new_n828_), .B2(new_n813_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n886_), .A2(new_n320_), .A3(new_n561_), .A4(new_n876_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n713_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n320_), .ZN(G1349gat));
  OR3_X1    g688(.A1(new_n886_), .A2(new_n603_), .A3(new_n876_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n603_), .A2(new_n411_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n890_), .A2(new_n317_), .B1(new_n883_), .B2(new_n891_), .ZN(G1350gat));
  NAND4_X1  g691(.A1(new_n883_), .A2(new_n410_), .A3(new_n409_), .A4(new_n619_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n883_), .A2(new_n533_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n291_), .ZN(G1351gat));
  NAND2_X1  g694(.A1(new_n861_), .A2(new_n875_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n582_), .ZN(new_n897_));
  INV_X1    g696(.A(G197gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1352gat));
  NOR2_X1   g698(.A1(new_n896_), .A2(new_n561_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT125), .B(G204gat), .Z(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n900_), .B2(new_n903_), .ZN(G1353gat));
  NOR2_X1   g703(.A1(new_n896_), .A2(new_n603_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n905_), .B2(new_n906_), .ZN(G1354gat));
  XOR2_X1   g708(.A(KEYINPUT126), .B(G218gat), .Z(new_n910_));
  NOR3_X1   g709(.A1(new_n896_), .A2(new_n653_), .A3(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n861_), .A2(new_n619_), .A3(new_n875_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n910_), .ZN(G1355gat));
endmodule


