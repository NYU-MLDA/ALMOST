//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT70), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT72), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(new_n203_), .B2(KEYINPUT35), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT8), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT65), .B(KEYINPUT66), .Z(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT7), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G85gat), .B(G92gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n209_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  AOI211_X1 g023(.A(KEYINPUT8), .B(new_n222_), .C1(new_n220_), .C2(new_n215_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT10), .B(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT9), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(G85gat), .A3(G92gat), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n215_), .B(new_n232_), .C1(new_n231_), .C2(new_n222_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n234_), .A2(KEYINPUT68), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(KEYINPUT68), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n226_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G29gat), .B(G36gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT15), .Z(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT71), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n237_), .A2(KEYINPUT71), .A3(new_n241_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n208_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n234_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n226_), .A2(new_n247_), .A3(KEYINPUT67), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n224_), .A2(new_n225_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n250_), .B2(new_n234_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(new_n240_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n206_), .B1(new_n246_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n246_), .A2(new_n206_), .A3(new_n254_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G190gat), .B(G218gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(G134gat), .B(G162gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(KEYINPUT36), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(KEYINPUT36), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n256_), .A2(new_n257_), .A3(new_n263_), .A4(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n257_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n262_), .B1(new_n266_), .B2(new_n255_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n265_), .A2(KEYINPUT37), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT37), .B1(new_n265_), .B2(new_n267_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271_));
  INV_X1    g070(.A(G1gat), .ZN(new_n272_));
  INV_X1    g071(.A(G8gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT14), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G1gat), .B(G8gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G231gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G57gat), .B(G64gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT11), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G71gat), .B(G78gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n282_), .A2(new_n283_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n280_), .A2(KEYINPUT11), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n279_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT17), .ZN(new_n291_));
  XOR2_X1   g090(.A(G127gat), .B(G155gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT16), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G183gat), .B(G211gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  OR3_X1    g094(.A1(new_n290_), .A2(new_n291_), .A3(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(KEYINPUT17), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n270_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT77), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT76), .B(KEYINPUT25), .ZN(new_n304_));
  INV_X1    g103(.A(G183gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT25), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n307_), .A2(KEYINPUT76), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(KEYINPUT76), .ZN(new_n309_));
  OAI211_X1 g108(.A(KEYINPUT77), .B(G183gat), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n312_), .A2(new_n313_), .B1(KEYINPUT25), .B2(new_n305_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n306_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(G169gat), .B2(G176gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT23), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G183gat), .A3(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NOR3_X1   g124(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n320_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n321_), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n324_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT78), .B1(new_n321_), .B2(KEYINPUT23), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n329_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G169gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT22), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT22), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G169gat), .ZN(new_n337_));
  INV_X1    g136(.A(G176gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n315_), .A2(new_n328_), .B1(new_n333_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT30), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345_));
  INV_X1    g144(.A(G43gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348_));
  INV_X1    g147(.A(G15gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n347_), .B(new_n350_), .Z(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n344_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n344_), .A2(new_n352_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT31), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G113gat), .B(G120gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n361_), .A2(KEYINPUT79), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n359_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(KEYINPUT79), .B2(new_n361_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT31), .B1(new_n353_), .B2(new_n354_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n357_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n357_), .B2(new_n366_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT19), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n373_));
  INV_X1    g172(.A(G218gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G211gat), .ZN(new_n375_));
  INV_X1    g174(.A(G211gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G218gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n379_));
  INV_X1    g178(.A(G204gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT21), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(G197gat), .B2(G204gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n378_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(G197gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n381_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n383_), .B(new_n386_), .C1(new_n387_), .C2(new_n380_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n387_), .B2(new_n380_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n383_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n385_), .A2(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n373_), .B1(new_n343_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n322_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(new_n330_), .A3(new_n324_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n312_), .A2(new_n313_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT25), .B(G183gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n326_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n395_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n339_), .A2(KEYINPUT89), .A3(new_n340_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n325_), .A2(new_n329_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT89), .B1(new_n339_), .B2(new_n340_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n400_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n385_), .A2(new_n388_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n389_), .A2(new_n390_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n372_), .B1(new_n392_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n372_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n315_), .A2(new_n328_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n342_), .A2(new_n333_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n391_), .A3(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n413_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n410_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT92), .ZN(new_n420_));
  XOR2_X1   g219(.A(G8gat), .B(G36gat), .Z(new_n421_));
  OR2_X1    g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n421_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n425_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n422_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n370_), .B1(new_n418_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n405_), .A2(new_n408_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n416_), .A3(KEYINPUT20), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n372_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n426_), .A2(new_n428_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n399_), .A2(new_n325_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n313_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n438_), .A2(new_n311_), .B1(new_n307_), .B2(G183gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(G183gat), .B1(new_n308_), .B2(new_n309_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n440_), .B2(new_n303_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n437_), .B1(new_n441_), .B2(new_n310_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n341_), .B1(new_n395_), .B2(new_n329_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n408_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n404_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(new_n391_), .A3(KEYINPUT90), .A4(new_n400_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n372_), .A2(new_n411_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n436_), .A2(new_n444_), .A3(new_n447_), .A4(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n433_), .A2(new_n434_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT97), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n433_), .A2(new_n434_), .A3(new_n449_), .A4(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n430_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  AND4_X1   g253(.A1(new_n436_), .A2(new_n444_), .A3(new_n447_), .A4(new_n448_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n413_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n429_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT27), .B1(new_n457_), .B2(new_n450_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT98), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n454_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n458_), .A2(new_n459_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT99), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n450_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n370_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT98), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT99), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n458_), .A2(new_n459_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .A4(new_n454_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n369_), .B1(new_n462_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT29), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G141gat), .A2(G148gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT82), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT2), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT2), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n472_), .A2(KEYINPUT82), .A3(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G141gat), .A2(G148gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT3), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n474_), .A2(new_n476_), .A3(new_n477_), .A4(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT83), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n477_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n486_), .A2(KEYINPUT83), .A3(new_n476_), .A4(new_n474_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G155gat), .A2(G162gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G155gat), .A2(G162gat), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n490_), .A2(KEYINPUT80), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(KEYINPUT80), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n489_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT84), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n488_), .A2(new_n497_), .A3(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n489_), .A2(KEYINPUT1), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n500_), .B(KEYINPUT81), .Z(new_n501_));
  OR2_X1    g300(.A1(new_n491_), .A2(new_n492_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n501_), .B(new_n502_), .C1(KEYINPUT1), .C2(new_n489_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n472_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(new_n478_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n471_), .B1(new_n499_), .B2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n497_), .B1(new_n488_), .B2(new_n494_), .ZN(new_n508_));
  AOI211_X1 g307(.A(KEYINPUT84), .B(new_n493_), .C1(new_n483_), .C2(new_n487_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n471_), .B(new_n506_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n470_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G22gat), .B(G50gat), .Z(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT85), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n510_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n470_), .A3(new_n513_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n515_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n513_), .B1(new_n519_), .B2(new_n470_), .ZN(new_n522_));
  AOI211_X1 g321(.A(KEYINPUT29), .B(new_n514_), .C1(new_n518_), .C2(new_n510_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT88), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n518_), .A2(KEYINPUT29), .A3(new_n510_), .ZN(new_n528_));
  AND2_X1   g327(.A1(G228gat), .A2(G233gat), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n391_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n496_), .A2(new_n498_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n408_), .B1(new_n532_), .B2(new_n470_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n529_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G78gat), .B(G106gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n531_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n527_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n531_), .A2(new_n534_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n535_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n531_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n526_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n525_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n539_), .A2(new_n543_), .B1(new_n524_), .B2(new_n521_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n469_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n521_), .A2(new_n524_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n537_), .A2(new_n538_), .A3(new_n527_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n526_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n525_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n460_), .A2(new_n461_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n550_), .A2(new_n369_), .A3(new_n551_), .A4(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n546_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n518_), .A2(new_n365_), .A3(new_n510_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n361_), .A2(new_n363_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n532_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G225gat), .A2(G233gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n555_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT95), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n555_), .A2(KEYINPUT4), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(KEYINPUT4), .A3(new_n557_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n558_), .B(KEYINPUT93), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G1gat), .B(G29gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT0), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G57gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT94), .B(G85gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  AND3_X1   g368(.A1(new_n560_), .A2(new_n564_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n554_), .A2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n574_), .A2(new_n456_), .A3(new_n455_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n418_), .B2(new_n574_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n570_), .A2(KEYINPUT33), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n560_), .A2(KEYINPUT33), .A3(new_n564_), .A4(new_n569_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n555_), .A2(new_n557_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n569_), .B1(new_n580_), .B2(new_n563_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n561_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n463_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n577_), .B1(new_n578_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n369_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n573_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n252_), .A2(new_n287_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n252_), .A2(new_n287_), .ZN(new_n592_));
  OAI211_X1 g391(.A(G230gat), .B(G233gat), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n252_), .B2(new_n287_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n237_), .A2(KEYINPUT12), .A3(new_n288_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n590_), .A4(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT5), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT69), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n593_), .A2(new_n598_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n603_), .B1(new_n593_), .B2(new_n598_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT13), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT13), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n277_), .A2(new_n240_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT73), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n241_), .A2(new_n277_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT74), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n615_), .A2(KEYINPUT74), .A3(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n277_), .A2(new_n240_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n613_), .A2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n622_), .A2(new_n616_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(G113gat), .B(G141gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT75), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G169gat), .B(G197gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n624_), .A2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n619_), .A2(new_n623_), .A3(new_n620_), .A4(new_n628_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n610_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n302_), .A2(new_n589_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n572_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n272_), .A3(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT38), .ZN(new_n639_));
  AOI22_X1  g438(.A1(new_n554_), .A2(new_n572_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n265_), .A2(new_n267_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n634_), .A3(new_n300_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT100), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(new_n637_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n639_), .B1(new_n646_), .B2(new_n272_), .ZN(G1324gat));
  NAND2_X1  g446(.A1(new_n462_), .A2(new_n468_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n636_), .A2(new_n273_), .A3(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n644_), .A2(new_n648_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT101), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n273_), .B1(new_n651_), .B2(KEYINPUT101), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n650_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  AOI21_X1  g458(.A(new_n349_), .B1(new_n645_), .B2(new_n586_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n661_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n636_), .A2(new_n349_), .A3(new_n586_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n544_), .A2(new_n545_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n645_), .B2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT42), .Z(new_n669_));
  NAND3_X1  g468(.A1(new_n636_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1327gat));
  NOR2_X1   g470(.A1(new_n641_), .A2(new_n300_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n589_), .A2(new_n634_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n637_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n676_), .B(new_n678_), .C1(new_n640_), .C2(new_n270_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  INV_X1    g479(.A(new_n270_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n589_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n585_), .A2(new_n587_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n637_), .B1(new_n546_), .B2(new_n553_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n676_), .B1(new_n686_), .B2(new_n678_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n634_), .B(new_n299_), .C1(new_n683_), .C2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n690_), .A2(G29gat), .A3(new_n637_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n689_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n675_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  OR2_X1    g492(.A1(new_n648_), .A2(G36gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n673_), .A2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n696_));
  XOR2_X1   g495(.A(new_n695_), .B(new_n696_), .Z(new_n697_));
  OR2_X1    g496(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n690_), .A2(new_n649_), .A3(new_n692_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G36gat), .ZN(new_n701_));
  NAND2_X1  g500(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n702_), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n704_), .B(new_n699_), .C1(new_n700_), .C2(G36gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1329gat));
  OAI21_X1  g505(.A(new_n346_), .B1(new_n673_), .B2(new_n369_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n690_), .A2(new_n692_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n586_), .A2(G43gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n674_), .B2(new_n667_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n690_), .A2(G50gat), .A3(new_n667_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n692_), .ZN(G1331gat));
  INV_X1    g513(.A(new_n610_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(new_n632_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n640_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n302_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT106), .Z(new_n720_));
  INV_X1    g519(.A(G57gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n637_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n643_), .A2(new_n300_), .A3(new_n716_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n572_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n726_), .A3(new_n649_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G64gat), .B1(new_n723_), .B2(new_n648_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT48), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n720_), .A2(new_n731_), .A3(new_n586_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G71gat), .B1(new_n723_), .B2(new_n369_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n720_), .A2(new_n737_), .A3(new_n667_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n667_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G78gat), .B1(new_n723_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(G1335gat));
  AOI21_X1  g542(.A(new_n270_), .B1(new_n573_), .B2(new_n588_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT103), .B1(new_n744_), .B2(new_n677_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n679_), .A3(new_n682_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n717_), .A2(new_n300_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n637_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G85gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n718_), .A2(new_n672_), .ZN(new_n751_));
  INV_X1    g550(.A(G85gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n637_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n751_), .B2(new_n753_), .ZN(G1336gat));
  NOR3_X1   g553(.A1(new_n751_), .A2(G92gat), .A3(new_n648_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n748_), .A2(new_n649_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G92gat), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT109), .Z(G1337gat));
  NOR3_X1   g557(.A1(new_n751_), .A2(new_n229_), .A3(new_n369_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n748_), .A2(new_n586_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G99gat), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT51), .Z(G1338gat));
  OR3_X1    g561(.A1(new_n751_), .A2(G106gat), .A3(new_n739_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n746_), .A2(KEYINPUT110), .A3(new_n667_), .A4(new_n747_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(G106gat), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n747_), .B(new_n667_), .C1(new_n683_), .C2(new_n687_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n764_), .B1(new_n766_), .B2(new_n769_), .ZN(new_n770_));
  AND4_X1   g569(.A1(new_n764_), .A2(new_n769_), .A3(G106gat), .A4(new_n765_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n763_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n763_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT119), .ZN(new_n777_));
  INV_X1    g576(.A(G113gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n632_), .A2(new_n604_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n595_), .A2(KEYINPUT55), .A3(new_n590_), .A4(new_n597_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(G230gat), .A4(G233gat), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n597_), .A2(new_n590_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(G230gat), .A3(G233gat), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n783_), .A2(KEYINPUT55), .A3(new_n595_), .A4(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n598_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n782_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n603_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n789_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n779_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n616_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n628_), .B1(new_n615_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n795_), .B2(new_n622_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n797_), .A2(KEYINPUT113), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(KEYINPUT113), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n631_), .A3(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n607_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n641_), .B1(new_n794_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT57), .B(new_n641_), .C1(new_n794_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n800_), .A2(new_n605_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n789_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n793_), .B1(new_n808_), .B2(KEYINPUT114), .ZN(new_n809_));
  INV_X1    g608(.A(new_n780_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n810_), .A2(new_n784_), .B1(new_n786_), .B2(new_n598_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n603_), .B1(new_n811_), .B2(new_n782_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(KEYINPUT56), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n807_), .B1(new_n809_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT58), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n813_), .B1(new_n812_), .B2(KEYINPUT56), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n808_), .A2(KEYINPUT114), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n793_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT115), .B1(new_n821_), .B2(new_n807_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n270_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n806_), .B1(new_n818_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT118), .B1(new_n825_), .B2(new_n300_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n818_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n806_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n299_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n610_), .A2(new_n632_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n834_));
  OR3_X1    g633(.A1(new_n833_), .A2(new_n301_), .A3(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n833_), .B2(new_n301_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n826_), .A2(new_n831_), .A3(new_n837_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n546_), .A2(new_n572_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(KEYINPUT117), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(KEYINPUT117), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n842_));
  NOR3_X1   g641(.A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n839_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n300_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n835_), .A2(new_n836_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n838_), .A2(new_n843_), .B1(KEYINPUT59), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n778_), .B1(new_n848_), .B2(new_n632_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n847_), .A2(G113gat), .A3(new_n633_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n777_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n838_), .A2(new_n843_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n847_), .A2(KEYINPUT59), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n632_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G113gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n850_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(KEYINPUT119), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n851_), .A2(new_n857_), .ZN(G1340gat));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n848_), .B2(new_n610_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n847_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n610_), .A2(new_n862_), .A3(new_n859_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n862_), .B2(new_n859_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n861_), .A2(new_n864_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n860_), .A2(new_n865_), .ZN(G1341gat));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n848_), .B2(new_n300_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n847_), .A2(G127gat), .A3(new_n299_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT120), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n852_), .A2(new_n300_), .A3(new_n853_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G127gat), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873_));
  INV_X1    g672(.A(new_n869_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n870_), .A2(new_n875_), .ZN(G1342gat));
  AOI21_X1  g675(.A(G134gat), .B1(new_n861_), .B2(new_n642_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n681_), .A2(G134gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT121), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n848_), .B2(new_n879_), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n845_), .A2(new_n846_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n667_), .A2(new_n369_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n572_), .A2(new_n649_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n632_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n610_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g689(.A1(new_n885_), .A2(new_n299_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT61), .B(G155gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n886_), .B2(new_n642_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n681_), .A2(G162gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT122), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n886_), .B2(new_n896_), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n637_), .A2(new_n648_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n586_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n667_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n837_), .B1(new_n845_), .B2(new_n830_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n825_), .A2(KEYINPUT118), .A3(new_n300_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n632_), .B(new_n900_), .C1(new_n901_), .C2(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(G169gat), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n903_), .B2(G169gat), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  AOI211_X1 g707(.A(KEYINPUT124), .B(new_n904_), .C1(new_n903_), .C2(G169gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n335_), .A2(new_n337_), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n908_), .A2(new_n909_), .B1(new_n910_), .B2(new_n903_), .ZN(G1348gat));
  AND2_X1   g710(.A1(new_n838_), .A2(new_n900_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G176gat), .B1(new_n912_), .B2(new_n610_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n881_), .A2(new_n667_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n899_), .A2(new_n338_), .A3(new_n715_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NAND4_X1  g715(.A1(new_n914_), .A2(new_n586_), .A3(new_n300_), .A4(new_n898_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n299_), .A2(new_n397_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n305_), .A2(new_n917_), .B1(new_n912_), .B2(new_n918_), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n912_), .A2(new_n642_), .A3(new_n396_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n838_), .A2(new_n681_), .A3(new_n900_), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n921_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT125), .B1(new_n921_), .B2(G190gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n920_), .B1(new_n922_), .B2(new_n923_), .ZN(G1351gat));
  NAND2_X1  g723(.A1(new_n883_), .A2(new_n898_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n632_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g727(.A1(new_n925_), .A2(new_n715_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n380_), .ZN(G1353gat));
  AOI21_X1  g729(.A(new_n299_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT126), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n883_), .A2(new_n898_), .A3(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n935_), .B2(new_n933_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n934_), .B1(new_n933_), .B2(new_n935_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n925_), .B2(new_n270_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n642_), .A2(new_n374_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n925_), .B2(new_n941_), .ZN(G1355gat));
endmodule


