//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT85), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G43gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT23), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OR3_X1    g012(.A1(new_n210_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT22), .B1(new_n210_), .B2(KEYINPUT84), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n211_), .A3(new_n215_), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n209_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n212_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT81), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT25), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT82), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(KEYINPUT82), .A3(new_n224_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n220_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n219_), .A2(new_n218_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n208_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT83), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n217_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n206_), .B(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G227gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(G15gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT86), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT30), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n239_), .B(new_n241_), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n234_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT87), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(G197gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT90), .B(G204gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(G197gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(G211gat), .B(G218gat), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n248_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT90), .B(G204gat), .Z(new_n254_));
  INV_X1    g053(.A(KEYINPUT91), .ZN(new_n255_));
  INV_X1    g054(.A(G197gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n245_), .A2(G197gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n255_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT21), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n249_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n261_), .A2(KEYINPUT92), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT92), .B1(new_n261_), .B2(new_n262_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n253_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(G228gat), .ZN(new_n266_));
  INV_X1    g065(.A(G233gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(KEYINPUT1), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(KEYINPUT1), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(KEYINPUT88), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(KEYINPUT88), .B2(new_n274_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  OR2_X1    g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT2), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n278_), .A2(KEYINPUT3), .B1(new_n280_), .B2(new_n277_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(KEYINPUT3), .B2(new_n278_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT89), .Z(new_n284_));
  OAI211_X1 g083(.A(new_n272_), .B(new_n271_), .C1(new_n282_), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n265_), .A2(new_n269_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n265_), .A2(KEYINPUT93), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT93), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n290_), .B(new_n253_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n287_), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n288_), .B1(new_n292_), .B2(new_n268_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G78gat), .B(G106gat), .Z(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT94), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT28), .B(G22gat), .ZN(new_n297_));
  INV_X1    g096(.A(G50gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n296_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT95), .B1(new_n295_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT95), .ZN(new_n303_));
  INV_X1    g102(.A(new_n294_), .ZN(new_n304_));
  AOI211_X1 g103(.A(new_n304_), .B(new_n288_), .C1(new_n292_), .C2(new_n268_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n303_), .B(new_n300_), .C1(new_n305_), .C2(KEYINPUT94), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n293_), .A2(new_n294_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(new_n305_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT97), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n204_), .B1(new_n286_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n204_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n279_), .A2(KEYINPUT97), .A3(new_n285_), .A4(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(KEYINPUT4), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n286_), .A2(new_n319_), .A3(new_n204_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n316_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n313_), .A2(new_n317_), .A3(new_n315_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G1gat), .B(G29gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT98), .B(G85gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT0), .B(G57gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n321_), .A2(new_n322_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n302_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT27), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT19), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n261_), .A2(new_n262_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT92), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n261_), .A2(KEYINPUT92), .A3(new_n262_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n252_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT20), .B1(new_n343_), .B2(new_n233_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT25), .B(G183gat), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n220_), .B1(new_n224_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n231_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT22), .B(G169gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n212_), .B1(new_n349_), .B2(new_n211_), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(KEYINPUT96), .Z(new_n351_));
  AOI21_X1  g150(.A(new_n348_), .B1(new_n351_), .B2(new_n209_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n352_), .B(new_n253_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n338_), .B1(new_n344_), .B2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n351_), .A2(new_n209_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n265_), .B1(new_n356_), .B2(new_n348_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n343_), .A2(new_n233_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT20), .A4(new_n337_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361_));
  INV_X1    g160(.A(G92gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT18), .B(G64gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n355_), .A2(new_n359_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n289_), .A2(new_n291_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n352_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n344_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n338_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AND4_X1   g172(.A1(KEYINPUT20), .A2(new_n357_), .A3(new_n338_), .A4(new_n358_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n367_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n335_), .B1(new_n360_), .B2(new_n365_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n335_), .A2(new_n369_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n311_), .A2(new_n333_), .A3(new_n334_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT100), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n379_), .B(KEYINPUT99), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n360_), .B2(new_n384_), .ZN(new_n385_));
  AOI211_X1 g184(.A(KEYINPUT100), .B(new_n383_), .C1(new_n355_), .C2(new_n359_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n381_), .B(new_n332_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n331_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n316_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n313_), .A2(new_n318_), .A3(new_n315_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n391_), .A2(new_n328_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n331_), .A2(new_n388_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n389_), .A2(new_n393_), .A3(new_n366_), .A4(new_n368_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n302_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n309_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n244_), .B1(new_n378_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n396_), .A2(new_n397_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n377_), .A2(new_n243_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n400_), .A2(new_n332_), .A3(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G230gat), .A2(G233gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G57gat), .A2(G64gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G57gat), .A2(G64gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT11), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT11), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n405_), .ZN(new_n411_));
  INV_X1    g210(.A(G71gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT66), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT66), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G71gat), .ZN(new_n415_));
  INV_X1    g214(.A(G78gat), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n408_), .B(new_n411_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(new_n415_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G78gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n410_), .B1(new_n409_), .B2(new_n405_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT67), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT67), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n419_), .A2(new_n427_), .A3(new_n424_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G85gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n362_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G85gat), .A2(G92gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT9), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT10), .B(G99gat), .Z(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n432_), .A2(KEYINPUT9), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n435_), .A2(new_n438_), .A3(new_n441_), .A4(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n444_));
  INV_X1    g243(.A(G99gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n437_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT64), .B1(new_n448_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n441_), .A2(new_n455_), .A3(new_n447_), .A4(new_n446_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n433_), .A2(KEYINPUT8), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT8), .ZN(new_n459_));
  INV_X1    g258(.A(new_n447_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n451_), .A2(KEYINPUT65), .A3(new_n452_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n459_), .B1(new_n466_), .B2(new_n434_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n443_), .B1(new_n458_), .B2(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT70), .B(new_n404_), .C1(new_n429_), .C2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT65), .B1(new_n451_), .B2(new_n452_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(new_n448_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n433_), .B1(new_n473_), .B2(new_n463_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n471_), .B1(new_n474_), .B2(new_n459_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n475_), .A2(new_n443_), .A3(new_n428_), .A4(new_n426_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT70), .B1(new_n476_), .B2(new_n404_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n470_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT69), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n419_), .A2(new_n479_), .A3(new_n424_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n481_), .A2(KEYINPUT12), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT68), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n475_), .B2(new_n443_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n484_), .B(new_n443_), .C1(new_n458_), .C2(new_n467_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n483_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT12), .B1(new_n429_), .B2(new_n468_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n429_), .A2(new_n468_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n492_), .A2(new_n476_), .ZN(new_n493_));
  OAI22_X1  g292(.A1(new_n478_), .A2(new_n491_), .B1(new_n493_), .B2(new_n404_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G176gat), .B(G204gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT72), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT71), .ZN(new_n497_));
  XOR2_X1   g296(.A(G120gat), .B(G148gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT5), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n497_), .B(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n494_), .A2(new_n500_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n503_), .A2(KEYINPUT13), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(KEYINPUT13), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT78), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT77), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT73), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G29gat), .B(G36gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n511_), .B(KEYINPUT73), .ZN(new_n516_));
  INV_X1    g315(.A(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520_));
  INV_X1    g319(.A(G1gat), .ZN(new_n521_));
  INV_X1    g320(.A(G8gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n519_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n515_), .A2(new_n518_), .A3(KEYINPUT15), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n510_), .B(new_n527_), .C1(new_n531_), .C2(new_n526_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n519_), .B(new_n526_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n510_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n509_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT77), .B1(new_n533_), .B2(new_n534_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n508_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G169gat), .B(G197gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT79), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n536_), .A2(new_n508_), .A3(new_n537_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT80), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n532_), .A2(new_n535_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n537_), .B1(new_n547_), .B2(KEYINPUT77), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT78), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT80), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n543_), .A4(new_n538_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n542_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n546_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n507_), .A2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n403_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n468_), .A2(KEYINPUT68), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n531_), .B1(new_n561_), .B2(new_n486_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT34), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT74), .B1(new_n565_), .B2(new_n566_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n519_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n570_), .B2(new_n468_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n562_), .A2(new_n568_), .A3(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n530_), .B(new_n529_), .C1(new_n485_), .C2(new_n487_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n571_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n567_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n560_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n568_), .B1(new_n562_), .B2(new_n571_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n567_), .A3(new_n574_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n560_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n558_), .A2(new_n559_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n577_), .B(new_n578_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT37), .B1(new_n582_), .B2(KEYINPUT75), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585_));
  AOI211_X1 g384(.A(new_n584_), .B(new_n585_), .C1(new_n576_), .C2(new_n581_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT76), .Z(new_n590_));
  XOR2_X1   g389(.A(new_n526_), .B(new_n590_), .Z(new_n591_));
  INV_X1    g390(.A(new_n482_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n591_), .A2(new_n592_), .A3(new_n480_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n480_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(G211gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT16), .B(G183gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  AND4_X1   g397(.A1(KEYINPUT17), .A2(new_n593_), .A3(new_n594_), .A4(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n591_), .B(new_n429_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n598_), .B(KEYINPUT17), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n588_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n555_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n555_), .A2(KEYINPUT101), .A3(new_n605_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n608_), .A2(new_n521_), .A3(new_n332_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n582_), .B(KEYINPUT102), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(new_n604_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n403_), .A2(new_n554_), .A3(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n333_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n610_), .A2(new_n611_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(new_n617_), .A3(new_n618_), .ZN(G1324gat));
  INV_X1    g418(.A(new_n377_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n608_), .A2(new_n522_), .A3(new_n620_), .A4(new_n609_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT103), .B1(new_n616_), .B2(new_n377_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(G8gat), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n616_), .A2(KEYINPUT103), .A3(new_n377_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n622_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  AND4_X1   g425(.A1(new_n622_), .A2(new_n625_), .A3(G8gat), .A4(new_n623_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n621_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT40), .B(new_n621_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1325gat));
  INV_X1    g431(.A(new_n244_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G15gat), .B1(new_n616_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT41), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(KEYINPUT41), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n608_), .A2(new_n609_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n244_), .A2(new_n236_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n635_), .B(new_n636_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(new_n400_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G22gat), .B1(new_n616_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT42), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n642_), .A2(G22gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n637_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(G1327gat));
  NOR2_X1   g447(.A1(new_n613_), .A2(new_n603_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n555_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(G29gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n332_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n588_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(new_n588_), .C1(new_n399_), .C2(new_n402_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n554_), .A2(new_n604_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT44), .B1(new_n658_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662_));
  AOI211_X1 g461(.A(new_n662_), .B(new_n659_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n661_), .A2(new_n663_), .A3(new_n333_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n653_), .B1(new_n664_), .B2(new_n652_), .ZN(G1328gat));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n666_), .A2(KEYINPUT107), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(KEYINPUT107), .ZN(new_n668_));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n661_), .A2(new_n663_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(new_n620_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n377_), .A2(G36gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n650_), .B2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n555_), .A2(new_n649_), .A3(new_n674_), .A4(new_n672_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n667_), .B(new_n668_), .C1(new_n671_), .C2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n661_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n658_), .A2(KEYINPUT44), .A3(new_n660_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n620_), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  INV_X1    g482(.A(new_n678_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n683_), .A2(KEYINPUT107), .A3(new_n666_), .A4(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n679_), .A2(new_n685_), .ZN(G1329gat));
  NAND3_X1  g485(.A1(new_n670_), .A2(G43gat), .A3(new_n243_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT108), .B(G43gat), .Z(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n650_), .B2(new_n633_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g491(.A1(new_n651_), .A2(new_n298_), .A3(new_n400_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n661_), .A2(new_n663_), .A3(new_n642_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT109), .ZN(new_n695_));
  OAI21_X1  g494(.A(G50gat), .B1(new_n694_), .B2(KEYINPUT109), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(G1331gat));
  INV_X1    g496(.A(new_n553_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n506_), .A2(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n403_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n615_), .ZN(new_n701_));
  INV_X1    g500(.A(G57gat), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n333_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n605_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n332_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n703_), .B1(new_n702_), .B2(new_n706_), .ZN(G1332gat));
  OAI21_X1  g506(.A(G64gat), .B1(new_n701_), .B2(new_n377_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT48), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n377_), .A2(G64gat), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT110), .Z(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n704_), .B2(new_n711_), .ZN(G1333gat));
  OAI21_X1  g511(.A(G71gat), .B1(new_n701_), .B2(new_n633_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT49), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT49), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(G71gat), .C1(new_n701_), .C2(new_n633_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n705_), .A2(new_n412_), .A3(new_n244_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n717_), .A2(KEYINPUT111), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1334gat));
  OAI21_X1  g522(.A(G78gat), .B1(new_n701_), .B2(new_n642_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n400_), .A2(new_n416_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT112), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n704_), .B2(new_n727_), .ZN(G1335gat));
  NAND2_X1  g527(.A1(new_n700_), .A2(new_n649_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G85gat), .B1(new_n730_), .B2(new_n332_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n699_), .A2(new_n604_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n658_), .A2(new_n733_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n734_), .A2(new_n430_), .A3(new_n333_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n731_), .A2(new_n735_), .ZN(G1336gat));
  AOI21_X1  g535(.A(G92gat), .B1(new_n730_), .B2(new_n620_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n734_), .A2(new_n362_), .A3(new_n377_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1337gat));
  INV_X1    g538(.A(new_n734_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n445_), .B1(new_n740_), .B2(new_n244_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n243_), .A2(new_n436_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n730_), .B2(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(G1338gat));
  NAND3_X1  g544(.A1(new_n730_), .A2(new_n437_), .A3(new_n400_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n658_), .A2(new_n400_), .A3(new_n733_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(G106gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n747_), .B2(G106gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g551(.A(G113gat), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n401_), .A2(new_n333_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n642_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n542_), .B1(new_n533_), .B2(new_n510_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n527_), .B1(new_n531_), .B2(new_n526_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n510_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n552_), .A2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(new_n502_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n481_), .A2(KEYINPUT12), .A3(new_n482_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n561_), .B2(new_n486_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n429_), .A2(new_n468_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n489_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n766_), .B2(new_n404_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n478_), .B2(new_n491_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n488_), .A2(new_n476_), .A3(new_n490_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n404_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(KEYINPUT115), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT70), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n765_), .B2(new_n771_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n469_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n764_), .A2(new_n489_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT55), .A3(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n767_), .A2(new_n769_), .A3(new_n772_), .A4(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n500_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n500_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT58), .B(new_n761_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n761_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n783_));
  AOI21_X1  g582(.A(new_n587_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n784_), .B2(KEYINPUT119), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT119), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n786_), .B(new_n587_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n779_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n778_), .A2(new_n500_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT116), .B(KEYINPUT56), .C1(new_n778_), .C2(new_n500_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n789_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n549_), .A2(new_n543_), .A3(new_n538_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n797_), .A2(KEYINPUT80), .B1(new_n548_), .B2(new_n542_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n502_), .B1(new_n798_), .B2(new_n551_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(new_n796_), .A3(new_n799_), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n503_), .A2(new_n760_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n796_), .B1(new_n795_), .B2(new_n799_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n613_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n788_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT57), .B(new_n613_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n603_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n506_), .A2(KEYINPUT114), .A3(new_n553_), .A4(new_n603_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n553_), .A2(new_n504_), .A3(new_n505_), .A4(new_n603_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n809_), .B1(new_n814_), .B2(new_n587_), .ZN(new_n815_));
  AOI211_X1 g614(.A(KEYINPUT54), .B(new_n588_), .C1(new_n810_), .C2(new_n813_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n756_), .B1(new_n808_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n753_), .B1(new_n818_), .B2(new_n553_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT120), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n753_), .C1(new_n818_), .C2(new_n553_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n818_), .B2(KEYINPUT59), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n804_), .A2(new_n805_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n788_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n807_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n817_), .B1(new_n829_), .B2(new_n604_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n824_), .B(KEYINPUT59), .C1(new_n830_), .C2(new_n755_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n830_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n756_), .A2(KEYINPUT122), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n756_), .A2(KEYINPUT122), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n833_), .A2(new_n834_), .A3(KEYINPUT59), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n826_), .A2(new_n831_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT123), .B(G113gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n553_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n823_), .B1(new_n836_), .B2(new_n838_), .ZN(G1340gat));
  NAND2_X1  g638(.A1(new_n832_), .A2(new_n835_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n831_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n507_), .B(new_n840_), .C1(new_n841_), .C2(new_n825_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G120gat), .ZN(new_n843_));
  INV_X1    g642(.A(new_n818_), .ZN(new_n844_));
  INV_X1    g643(.A(G120gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n506_), .B2(KEYINPUT60), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n844_), .B(new_n846_), .C1(KEYINPUT60), .C2(new_n845_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n847_), .ZN(G1341gat));
  AOI21_X1  g647(.A(G127gat), .B1(new_n844_), .B2(new_n603_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n603_), .A2(G127gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n836_), .B2(new_n850_), .ZN(G1342gat));
  AOI21_X1  g650(.A(G134gat), .B1(new_n844_), .B2(new_n614_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n588_), .A2(G134gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n836_), .B2(new_n853_), .ZN(G1343gat));
  NOR4_X1   g653(.A1(new_n642_), .A2(new_n333_), .A3(new_n620_), .A4(new_n244_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n832_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n698_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n507_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  OAI211_X1 g659(.A(new_n603_), .B(new_n855_), .C1(new_n808_), .C2(new_n817_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n861_), .A2(KEYINPUT124), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(KEYINPUT124), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1346gat));
  AOI21_X1  g666(.A(G162gat), .B1(new_n856_), .B2(new_n614_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n588_), .A2(G162gat), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n856_), .B2(new_n869_), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n830_), .A2(new_n377_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n633_), .A2(new_n400_), .A3(new_n332_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873_), .B2(new_n553_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT62), .B(G169gat), .C1(new_n873_), .C2(new_n553_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n871_), .A2(new_n698_), .A3(new_n349_), .A4(new_n872_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(G1348gat));
  NOR2_X1   g678(.A1(new_n873_), .A2(new_n506_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n211_), .ZN(G1349gat));
  NOR2_X1   g680(.A1(new_n873_), .A2(new_n604_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n345_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n221_), .B2(new_n882_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n873_), .B2(new_n587_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n614_), .A2(new_n224_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n873_), .B2(new_n886_), .ZN(G1351gat));
  NAND2_X1  g686(.A1(new_n400_), .A2(new_n333_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n244_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n620_), .B(new_n889_), .C1(new_n808_), .C2(new_n817_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n891_), .A2(new_n698_), .B1(KEYINPUT125), .B2(G197gat), .ZN(new_n892_));
  OR2_X1    g691(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1352gat));
  NOR2_X1   g693(.A1(new_n890_), .A2(new_n506_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n247_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n245_), .B2(new_n895_), .ZN(G1353gat));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT63), .B(G211gat), .Z(new_n899_));
  NAND4_X1  g698(.A1(new_n891_), .A2(new_n898_), .A3(new_n603_), .A4(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n891_), .A2(new_n603_), .A3(new_n899_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(KEYINPUT126), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n890_), .B2(new_n604_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT127), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n906_), .B(new_n903_), .C1(new_n890_), .C2(new_n604_), .ZN(new_n907_));
  AND4_X1   g706(.A1(new_n900_), .A2(new_n902_), .A3(new_n905_), .A4(new_n907_), .ZN(G1354gat));
  INV_X1    g707(.A(G218gat), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n890_), .A2(new_n909_), .A3(new_n587_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n891_), .A2(new_n614_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n909_), .ZN(G1355gat));
endmodule


