//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT114), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(KEYINPUT11), .B2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT67), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n206_), .B(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n208_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT12), .B1(new_n209_), .B2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT6), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  OR3_X1    g022(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT9), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n217_), .A2(new_n219_), .A3(new_n221_), .A4(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT69), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OR3_X1    g028(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n228_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n221_), .A2(new_n229_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n218_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT66), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n218_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT8), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n232_), .A2(new_n238_), .A3(new_n218_), .A4(new_n233_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n226_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n235_), .A2(new_n237_), .A3(KEYINPUT68), .A4(new_n239_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n214_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n209_), .A2(new_n213_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n240_), .A2(new_n225_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT12), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n244_), .A2(new_n245_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(new_n243_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n214_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT70), .ZN(new_n254_));
  AND2_X1   g053(.A1(G230gat), .A2(G233gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n247_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n209_), .A2(new_n213_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n257_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n248_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n255_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G120gat), .B(G148gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n259_), .A2(new_n262_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT13), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(KEYINPUT13), .A3(new_n271_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G8gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT79), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n278_), .A2(new_n279_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G15gat), .B(G22gat), .Z(new_n282_));
  NOR3_X1   g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G1gat), .B(G8gat), .Z(new_n284_));
  OR2_X1    g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n284_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G29gat), .B(G36gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G43gat), .B(G50gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT15), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n285_), .A2(new_n286_), .A3(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G229gat), .A2(G233gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n287_), .B(new_n290_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(new_n294_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G113gat), .B(G141gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT83), .ZN(new_n299_));
  XOR2_X1   g098(.A(G169gat), .B(G197gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n297_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n203_), .B1(new_n276_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G231gat), .A2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n287_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(new_n246_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT81), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G127gat), .B(G155gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(G183gat), .B(G211gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT17), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT82), .Z(new_n317_));
  NAND3_X1  g116(.A1(new_n309_), .A2(new_n310_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n315_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n307_), .A2(KEYINPUT17), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n274_), .A2(KEYINPUT114), .A3(new_n302_), .A4(new_n275_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n304_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT115), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT27), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT19), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n331_));
  INV_X1    g130(.A(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(G176gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT22), .B(G169gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n333_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n336_), .A2(KEYINPUT102), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT85), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(KEYINPUT85), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT23), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(G183gat), .B2(G190gat), .ZN(new_n343_));
  OAI22_X1  g142(.A1(new_n341_), .A2(new_n343_), .B1(G183gat), .B2(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n336_), .A2(KEYINPUT102), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n337_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n339_), .A2(new_n340_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(KEYINPUT23), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT100), .B(KEYINPUT24), .Z(new_n351_));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT101), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT101), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n350_), .A2(new_n357_), .A3(new_n354_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G169gat), .B(G176gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(G190gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT25), .B(G183gat), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n361_), .A2(new_n351_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n347_), .B1(new_n359_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT97), .ZN(new_n366_));
  INV_X1    g165(.A(G211gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n367_), .A2(G218gat), .ZN(new_n368_));
  INV_X1    g167(.A(G218gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n369_), .A2(G211gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n366_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(G211gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(G218gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(KEYINPUT97), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT99), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT99), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n371_), .A2(new_n377_), .A3(new_n374_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT95), .ZN(new_n379_));
  INV_X1    g178(.A(G197gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(G204gat), .ZN(new_n381_));
  INV_X1    g180(.A(G204gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n381_), .A2(new_n383_), .B1(new_n380_), .B2(G204gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT21), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n376_), .A2(new_n378_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT94), .B1(new_n382_), .B2(G197gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT93), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n380_), .B2(G204gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT94), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(new_n380_), .A3(G204gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n382_), .A2(KEYINPUT93), .A3(G197gat), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n389_), .A2(new_n391_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(KEYINPUT21), .A2(new_n395_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n380_), .A2(G204gat), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n382_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT95), .B1(new_n382_), .B2(G197gat), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n385_), .B(new_n397_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT96), .B1(new_n384_), .B2(new_n385_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n396_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT98), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n401_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n384_), .A2(KEYINPUT96), .A3(new_n385_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT98), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n396_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n388_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n331_), .B1(new_n365_), .B2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(KEYINPUT84), .B(G183gat), .Z(new_n413_));
  INV_X1    g212(.A(KEYINPUT25), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n362_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n343_), .B1(new_n349_), .B2(new_n342_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT24), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n352_), .A2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(new_n360_), .B2(new_n419_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n413_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n350_), .A2(new_n424_), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n335_), .A2(KEYINPUT86), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n332_), .A2(KEYINPUT22), .ZN(new_n427_));
  AOI21_X1  g226(.A(G176gat), .B1(new_n427_), .B2(KEYINPUT86), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n334_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n417_), .A2(new_n422_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n411_), .A2(KEYINPUT103), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT103), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n408_), .A2(new_n409_), .A3(new_n396_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n409_), .B1(new_n408_), .B2(new_n396_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n387_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n430_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n432_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n330_), .B(new_n412_), .C1(new_n431_), .C2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G8gat), .B(G36gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT104), .B(KEYINPUT18), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n430_), .B(new_n387_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(KEYINPUT20), .C1(new_n365_), .C2(new_n411_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n329_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n438_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n444_), .B1(new_n438_), .B2(new_n447_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n327_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT111), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT111), .B(new_n327_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G141gat), .ZN(new_n455_));
  INV_X1    g254(.A(G148gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G141gat), .A2(G148gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT91), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G155gat), .A2(G162gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT1), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n457_), .B(new_n458_), .C1(new_n461_), .C2(new_n463_), .ZN(new_n464_));
  OR3_X1    g263(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT2), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n458_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n465_), .A2(new_n467_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n459_), .B(KEYINPUT91), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n462_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n464_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT29), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n411_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G78gat), .B(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G228gat), .A2(G233gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT92), .B1(new_n477_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n480_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(new_n411_), .B2(new_n476_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n474_), .A2(new_n475_), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n485_), .B(KEYINPUT28), .Z(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G22gat), .B(G50gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(new_n491_), .A3(new_n489_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n448_), .A2(new_n327_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n446_), .A2(new_n329_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(KEYINPUT110), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n446_), .A2(new_n329_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n358_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n357_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n364_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n346_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT20), .B1(new_n503_), .B2(new_n435_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT103), .B1(new_n411_), .B2(new_n430_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n435_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n499_), .B1(new_n507_), .B2(new_n330_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n498_), .B1(new_n508_), .B2(KEYINPUT110), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n496_), .B1(new_n509_), .B2(new_n444_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G71gat), .B(G99gat), .ZN(new_n511_));
  INV_X1    g310(.A(G43gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT30), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n430_), .B(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT87), .B(G15gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G134gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G127gat), .ZN(new_n519_));
  INV_X1    g318(.A(G127gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G134gat), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT89), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(KEYINPUT89), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G113gat), .B(G120gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n524_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(new_n522_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT31), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT88), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G227gat), .A2(G233gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  OR2_X1    g333(.A1(new_n517_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n517_), .A2(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n473_), .A2(new_n530_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n464_), .A2(new_n526_), .A3(new_n472_), .A4(new_n529_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G225gat), .A2(G233gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(KEYINPUT105), .Z(new_n542_));
  NOR2_X1   g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n538_), .A2(KEYINPUT4), .A3(new_n539_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n473_), .A2(new_n530_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT106), .B(KEYINPUT0), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT107), .ZN(new_n551_));
  XOR2_X1   g350(.A(G1gat), .B(G29gat), .Z(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  XNOR2_X1  g352(.A(G57gat), .B(G85gat), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n554_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n549_), .B(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n537_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n454_), .A2(new_n495_), .A3(new_n510_), .A4(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT112), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n505_), .A2(new_n506_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n330_), .B1(new_n562_), .B2(new_n412_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT110), .B1(new_n563_), .B2(new_n497_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n498_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n443_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n452_), .A2(new_n453_), .B1(new_n567_), .B2(new_n496_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT112), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n495_), .A4(new_n559_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n558_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n438_), .A2(new_n447_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n443_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n438_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT111), .B1(new_n575_), .B2(new_n327_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n453_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n571_), .B(new_n510_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n555_), .A2(new_n556_), .B1(new_n542_), .B2(new_n540_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n545_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n580_), .A2(KEYINPUT108), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(KEYINPUT108), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT33), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n549_), .A2(new_n557_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n549_), .A2(KEYINPUT33), .A3(new_n557_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n586_), .A2(new_n573_), .A3(new_n574_), .A4(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT109), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n444_), .A2(KEYINPUT32), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n572_), .B2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n438_), .A2(KEYINPUT109), .A3(new_n447_), .A4(new_n590_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n558_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n590_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n588_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n495_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n578_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n537_), .B(KEYINPUT90), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n561_), .A2(new_n570_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n251_), .A2(new_n291_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT72), .ZN(new_n602_));
  INV_X1    g401(.A(new_n291_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT72), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n240_), .A2(new_n290_), .A3(new_n225_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT34), .Z(new_n609_));
  INV_X1    g408(.A(KEYINPUT35), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT73), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(KEYINPUT73), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n602_), .A2(new_n606_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n609_), .A2(new_n610_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT75), .ZN(new_n617_));
  INV_X1    g416(.A(new_n612_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n616_), .B(KEYINPUT74), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n617_), .B1(new_n620_), .B2(new_n604_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n601_), .A2(KEYINPUT75), .A3(new_n618_), .A4(new_n619_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n615_), .A2(new_n616_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT36), .Z(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n615_), .A2(new_n616_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n621_), .A2(new_n622_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n600_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n326_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n202_), .B1(new_n637_), .B2(new_n558_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n633_), .B(new_n640_), .C1(new_n623_), .C2(new_n628_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT78), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT78), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n629_), .A2(new_n643_), .A3(new_n640_), .A4(new_n633_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n627_), .B(KEYINPUT76), .Z(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT77), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT77), .B1(new_n623_), .B2(new_n646_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n633_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT37), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n321_), .B1(new_n645_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR4_X1   g453(.A1(new_n654_), .A2(new_n600_), .A3(new_n303_), .A4(new_n276_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n202_), .A3(new_n558_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n638_), .B1(new_n639_), .B2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n639_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(KEYINPUT113), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(KEYINPUT113), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(new_n568_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n655_), .A2(new_n277_), .A3(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n326_), .A2(new_n662_), .A3(new_n636_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(G8gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n664_), .B2(G8gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT40), .B(new_n663_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  INV_X1    g471(.A(G15gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n599_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n655_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n326_), .A2(new_n674_), .A3(new_n636_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n676_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT41), .B1(new_n676_), .B2(G15gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT116), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT116), .B(new_n675_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1326gat));
  INV_X1    g482(.A(G22gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n495_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n655_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n637_), .A2(new_n685_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G22gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT117), .B(KEYINPUT42), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n688_), .A2(new_n689_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n686_), .B1(new_n690_), .B2(new_n691_), .ZN(G1327gat));
  AND2_X1   g491(.A1(new_n304_), .A2(new_n323_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n321_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n561_), .A2(new_n570_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n598_), .A2(new_n599_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  AOI22_X1  g497(.A1(new_n644_), .A2(new_n642_), .B1(new_n651_), .B2(KEYINPUT37), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n645_), .A2(new_n652_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n600_), .B2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n694_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT118), .B(KEYINPUT44), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n693_), .A2(new_n321_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n698_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n600_), .A2(KEYINPUT43), .A3(new_n701_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n706_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n705_), .A2(G29gat), .A3(new_n558_), .A4(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n600_), .A2(new_n303_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n635_), .A2(new_n321_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n276_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G29gat), .B1(new_n716_), .B2(new_n558_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n711_), .A2(new_n717_), .ZN(G1328gat));
  OAI211_X1 g517(.A(new_n709_), .B(new_n662_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G36gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n568_), .A2(G36gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n712_), .A2(new_n714_), .A3(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT45), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(KEYINPUT46), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1329gat));
  NOR2_X1   g527(.A1(new_n537_), .A2(new_n512_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n709_), .B(new_n729_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n512_), .B1(new_n715_), .B2(new_n599_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g532(.A1(new_n705_), .A2(G50gat), .A3(new_n685_), .A4(new_n709_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G50gat), .B1(new_n716_), .B2(new_n685_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1331gat));
  INV_X1    g536(.A(new_n276_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(new_n302_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n636_), .A2(new_n322_), .A3(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(G57gat), .A3(new_n558_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT119), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(KEYINPUT119), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n697_), .A2(new_n739_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(new_n654_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G57gat), .B1(new_n745_), .B2(new_n558_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n742_), .A2(new_n743_), .A3(new_n746_), .ZN(G1332gat));
  INV_X1    g546(.A(G64gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n740_), .B2(new_n662_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT48), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(new_n748_), .A3(new_n662_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n740_), .B2(new_n674_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT49), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n745_), .A2(new_n753_), .A3(new_n674_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1334gat));
  INV_X1    g556(.A(G78gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n740_), .B2(new_n685_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT50), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n745_), .A2(new_n758_), .A3(new_n685_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1335gat));
  NOR2_X1   g561(.A1(new_n744_), .A2(new_n713_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n222_), .A3(new_n558_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n707_), .A2(new_n708_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n558_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n738_), .A2(new_n302_), .A3(new_n322_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n765_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n769_), .B2(new_n222_), .ZN(G1336gat));
  NAND3_X1  g569(.A1(new_n763_), .A2(new_n223_), .A3(new_n662_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n765_), .A2(new_n568_), .A3(new_n768_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n223_), .ZN(G1337gat));
  NOR3_X1   g572(.A1(new_n765_), .A2(new_n599_), .A3(new_n768_), .ZN(new_n774_));
  INV_X1    g573(.A(G99gat), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n763_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n535_), .A2(new_n536_), .A3(new_n215_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT51), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781_));
  OAI221_X1 g580(.A(new_n781_), .B1(new_n777_), .B2(new_n778_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n763_), .A2(new_n216_), .A3(new_n685_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n685_), .B(new_n767_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n784_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  OR2_X1    g592(.A1(new_n297_), .A2(new_n301_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n294_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n292_), .A2(new_n293_), .A3(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n301_), .C1(new_n296_), .C2(new_n795_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n271_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n251_), .A2(new_n252_), .A3(new_n245_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n248_), .A2(new_n249_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n244_), .A2(new_n245_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n804_), .A2(KEYINPUT120), .A3(KEYINPUT55), .A4(new_n258_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n250_), .A2(new_n254_), .A3(KEYINPUT55), .A4(new_n258_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n259_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n250_), .A2(new_n260_), .A3(new_n254_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n255_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n805_), .A2(new_n808_), .A3(new_n810_), .A4(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n268_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n799_), .B1(new_n814_), .B2(KEYINPUT56), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n816_), .A3(new_n268_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(KEYINPUT58), .A3(new_n817_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n699_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(KEYINPUT122), .A2(KEYINPUT57), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n816_), .A2(KEYINPUT121), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n814_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n813_), .A2(KEYINPUT121), .A3(new_n816_), .A4(new_n268_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n271_), .A2(new_n302_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n826_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n272_), .A2(new_n798_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n634_), .B(new_n824_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n828_), .B1(new_n814_), .B2(new_n825_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n831_), .B1(new_n833_), .B2(new_n827_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n823_), .B1(new_n834_), .B2(new_n635_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n822_), .A2(new_n832_), .A3(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n701_), .A2(new_n303_), .A3(new_n322_), .A4(new_n738_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT54), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n653_), .A2(new_n839_), .A3(new_n303_), .A4(new_n738_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n836_), .A2(new_n321_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  OR4_X1    g640(.A1(new_n537_), .A2(new_n662_), .A3(new_n766_), .A4(new_n685_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n302_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n836_), .A2(new_n321_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n838_), .A2(new_n840_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n842_), .A2(KEYINPUT123), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n842_), .A2(KEYINPUT123), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .A4(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n842_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n852_), .A2(new_n302_), .A3(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n845_), .B1(new_n854_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n738_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n843_), .B(new_n857_), .C1(KEYINPUT60), .C2(new_n856_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n852_), .A2(new_n276_), .A3(new_n853_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n856_), .ZN(G1341gat));
  NAND3_X1  g659(.A1(new_n843_), .A2(new_n520_), .A3(new_n322_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n852_), .A2(new_n322_), .A3(new_n853_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n520_), .ZN(G1342gat));
  NAND3_X1  g662(.A1(new_n843_), .A2(new_n518_), .A3(new_n635_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n852_), .A2(new_n699_), .A3(new_n853_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n518_), .ZN(G1343gat));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n568_), .A2(new_n599_), .A3(new_n558_), .A4(new_n685_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n848_), .B2(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n841_), .A2(KEYINPUT124), .A3(new_n868_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n302_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G141gat), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n455_), .B(new_n302_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1344gat));
  OAI21_X1  g674(.A(new_n276_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G148gat), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n456_), .B(new_n276_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1345gat));
  OAI21_X1  g678(.A(new_n322_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n881_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n322_), .B(new_n883_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1346gat));
  INV_X1    g684(.A(G162gat), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n886_), .B(new_n635_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n848_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT124), .B1(new_n841_), .B2(new_n868_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n701_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n886_), .B2(new_n890_), .ZN(G1347gat));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n568_), .A2(new_n599_), .A3(new_n558_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT125), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n894_), .A2(new_n685_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n848_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n303_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n892_), .B1(new_n898_), .B2(new_n332_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n335_), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT62), .B(G169gat), .C1(new_n897_), .C2(new_n303_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(G1348gat));
  AOI21_X1  g701(.A(new_n895_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n276_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g704(.A(new_n413_), .B1(new_n903_), .B2(new_n322_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n363_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n841_), .A2(new_n907_), .A3(new_n321_), .A4(new_n895_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT126), .B1(new_n906_), .B2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n903_), .A2(new_n363_), .A3(new_n322_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n841_), .A2(new_n321_), .A3(new_n895_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n910_), .B(new_n911_), .C1(new_n413_), .C2(new_n912_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n909_), .A2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n897_), .B2(new_n701_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n903_), .A2(new_n362_), .A3(new_n635_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1351gat));
  AND3_X1   g716(.A1(new_n662_), .A2(new_n599_), .A3(new_n571_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n848_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n303_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n380_), .ZN(G1352gat));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n738_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n382_), .ZN(G1353gat));
  INV_X1    g722(.A(new_n919_), .ZN(new_n924_));
  AND2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  AOI211_X1 g725(.A(new_n925_), .B(new_n321_), .C1(KEYINPUT127), .C2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n924_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(KEYINPUT127), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n924_), .B(new_n927_), .C1(KEYINPUT127), .C2(new_n926_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1354gat));
  OAI21_X1  g731(.A(G218gat), .B1(new_n919_), .B2(new_n701_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n635_), .A2(new_n369_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n919_), .B2(new_n934_), .ZN(G1355gat));
endmodule


