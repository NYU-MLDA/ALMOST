//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT86), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n205_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT87), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n205_), .A3(new_n209_), .ZN(new_n213_));
  AND3_X1   g012(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT87), .ZN(new_n217_));
  INV_X1    g016(.A(new_n211_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(new_n213_), .A3(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228_));
  NOR4_X1   g027(.A1(new_n228_), .A2(KEYINPUT88), .A3(G141gat), .A4(G148gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT88), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT3), .B1(new_n221_), .B2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n227_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(KEYINPUT89), .B(new_n227_), .C1(new_n229_), .C2(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n218_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT90), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT90), .ZN(new_n240_));
  AOI211_X1 g039(.A(new_n240_), .B(new_n237_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n204_), .B(new_n224_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n221_), .A2(new_n230_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n228_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n221_), .A2(new_n230_), .A3(KEYINPUT3), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT89), .B1(new_n247_), .B2(new_n227_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n235_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n238_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n240_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n236_), .A2(KEYINPUT90), .A3(new_n238_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n243_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n204_), .B(KEYINPUT85), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n242_), .B(KEYINPUT4), .C1(new_n253_), .C2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n224_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT97), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n256_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(new_n254_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(new_n242_), .A3(new_n260_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G29gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G85gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT0), .B(G57gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n263_), .A2(new_n265_), .A3(new_n270_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(KEYINPUT99), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT99), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n266_), .A2(new_n275_), .A3(new_n271_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT100), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(KEYINPUT100), .A3(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT31), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n254_), .B(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(KEYINPUT82), .A2(G183gat), .A3(G190gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT82), .B1(G183gat), .B2(G190gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT23), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT83), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n289_));
  INV_X1    g088(.A(G183gat), .ZN(new_n290_));
  INV_X1    g089(.A(G190gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT83), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n294_), .B(KEYINPUT23), .C1(new_n285_), .C2(new_n286_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n288_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT80), .B(G190gat), .Z(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(G183gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT84), .ZN(new_n300_));
  INV_X1    g099(.A(G169gat), .ZN(new_n301_));
  INV_X1    g100(.A(G176gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT22), .B(G169gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(new_n302_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n296_), .A2(new_n306_), .A3(new_n298_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n300_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n285_), .A2(new_n286_), .ZN(new_n309_));
  OAI22_X1  g108(.A1(new_n309_), .A2(KEYINPUT23), .B1(new_n292_), .B2(new_n289_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT24), .B1(new_n301_), .B2(new_n302_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  MUX2_X1   g111(.A(new_n311_), .B(KEYINPUT24), .S(new_n312_), .Z(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT25), .B(G183gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT26), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G190gat), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n314_), .B(new_n316_), .C1(new_n297_), .C2(new_n315_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n308_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n284_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G71gat), .B(G99gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G43gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT30), .B(G15gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n324_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n257_), .A2(KEYINPUT29), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT94), .ZN(new_n330_));
  INV_X1    g129(.A(G197gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(G204gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT21), .B(new_n332_), .C1(new_n334_), .C2(new_n330_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G211gat), .B(G218gat), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n334_), .A2(KEYINPUT95), .A3(KEYINPUT21), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT95), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT21), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n333_), .B2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n335_), .B(new_n336_), .C1(new_n337_), .C2(new_n340_), .ZN(new_n341_));
  OR3_X1    g140(.A1(new_n333_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n329_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G228gat), .ZN(new_n348_));
  INV_X1    g147(.A(G233gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n329_), .A2(new_n352_), .A3(new_n346_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G78gat), .B(G106gat), .Z(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n354_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n352_), .B1(new_n329_), .B2(new_n346_), .ZN(new_n357_));
  AOI211_X1 g156(.A(new_n350_), .B(new_n345_), .C1(new_n257_), .C2(KEYINPUT29), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G22gat), .B(G50gat), .Z(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n257_), .B2(KEYINPUT29), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  INV_X1    g162(.A(new_n361_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n253_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT92), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(new_n365_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT92), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n360_), .A2(new_n369_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT96), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n355_), .B2(new_n359_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n354_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n379_));
  OAI22_X1  g178(.A1(new_n379_), .A2(KEYINPUT96), .B1(new_n367_), .B2(new_n368_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n376_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383_));
  INV_X1    g182(.A(G92gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT18), .B(G64gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n319_), .B2(new_n343_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n343_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n310_), .B1(G183gat), .B2(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n305_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n291_), .A2(KEYINPUT26), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n316_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n314_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n296_), .A2(new_n313_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n390_), .A2(new_n392_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n389_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT19), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n308_), .A2(new_n390_), .A3(new_n318_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n392_), .A2(new_n397_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n388_), .B1(new_n405_), .B2(new_n343_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(new_n402_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n387_), .B1(new_n403_), .B2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n401_), .B1(new_n389_), .B2(new_n398_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n387_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n411_), .A2(new_n408_), .A3(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n382_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n411_), .B2(new_n408_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT98), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n405_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n392_), .A2(KEYINPUT98), .A3(new_n397_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n390_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n402_), .B1(new_n389_), .B2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n407_), .A2(new_n401_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n415_), .B(KEYINPUT27), .C1(new_n422_), .C2(new_n412_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n414_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n381_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n281_), .A2(new_n328_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n412_), .A2(KEYINPUT32), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n422_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n427_), .B1(new_n411_), .B2(new_n408_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n274_), .A2(new_n428_), .A3(new_n276_), .A4(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n410_), .A2(new_n413_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n273_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n256_), .A2(new_n260_), .A3(new_n259_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n264_), .A2(new_n242_), .A3(new_n262_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n271_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n273_), .A2(new_n432_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n431_), .A2(new_n433_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n381_), .B1(new_n430_), .B2(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n369_), .A2(new_n375_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n357_), .A2(new_n358_), .A3(new_n356_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT96), .B1(new_n379_), .B2(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n359_), .A2(new_n377_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n440_), .A2(new_n360_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n414_), .A2(new_n423_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n439_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n426_), .B1(new_n447_), .B2(new_n328_), .ZN(new_n448_));
  INV_X1    g247(.A(G1gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT74), .B(G8gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT14), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G15gat), .B(G22gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n449_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT14), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n452_), .A2(new_n454_), .A3(new_n449_), .ZN(new_n455_));
  OR3_X1    g254(.A1(new_n453_), .A2(new_n455_), .A3(G8gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(G8gat), .B1(new_n453_), .B2(new_n455_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G231gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G57gat), .ZN(new_n461_));
  INV_X1    g260(.A(G64gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT11), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G57gat), .A2(G64gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n467_));
  INV_X1    g266(.A(G78gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G71gat), .ZN(new_n469_));
  INV_X1    g268(.A(G71gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G78gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n467_), .B1(new_n466_), .B2(new_n472_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n464_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(G57gat), .A2(G64gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(G57gat), .A2(G64gat), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT11), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G71gat), .B(G78gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT67), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n466_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n475_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n477_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT75), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n460_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G127gat), .B(G155gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G211gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT16), .B(G183gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(new_n488_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT68), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n477_), .B2(new_n484_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n476_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n482_), .A2(new_n483_), .A3(new_n475_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(KEYINPUT68), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n460_), .B(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n492_), .B(KEYINPUT17), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n493_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT65), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT64), .ZN(new_n506_));
  INV_X1    g305(.A(G85gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(G92gat), .A3(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n507_), .A2(new_n384_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n510_), .A2(new_n511_), .B1(KEYINPUT9), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT6), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT10), .B(G99gat), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n516_), .B(new_n517_), .C1(new_n518_), .C2(G106gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n505_), .B1(new_n513_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n512_), .A2(KEYINPUT9), .ZN(new_n521_));
  AND2_X1   g320(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n384_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n511_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n521_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G99gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT10), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT10), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(G99gat), .ZN(new_n530_));
  AOI21_X1  g329(.A(G106gat), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n516_), .A2(new_n517_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n526_), .A2(KEYINPUT65), .A3(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n520_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G29gat), .B(G36gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G85gat), .B(G92gat), .Z(new_n539_));
  OR2_X1    g338(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n516_), .A2(new_n540_), .A3(new_n517_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n542_));
  INV_X1    g341(.A(G106gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n527_), .A3(new_n543_), .ZN(new_n544_));
  OAI211_X1 g343(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n539_), .B1(new_n541_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT8), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT8), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n549_), .B(new_n539_), .C1(new_n541_), .C2(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n535_), .A2(new_n538_), .A3(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n553_));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n552_), .B1(KEYINPUT35), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n538_), .B(KEYINPUT15), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n520_), .A2(new_n534_), .A3(KEYINPUT69), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT69), .B1(new_n520_), .B2(new_n534_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n551_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n556_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(KEYINPUT35), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n563_), .A2(KEYINPUT36), .A3(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n566_), .B(KEYINPUT36), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT37), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n568_), .A2(new_n573_), .A3(new_n570_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n504_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT72), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n551_), .A2(new_n534_), .A3(new_n520_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n499_), .A2(new_n579_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n495_), .A2(new_n498_), .B1(new_n535_), .B2(new_n551_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n578_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT5), .B(G176gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT71), .B(G204gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G120gat), .B(G148gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT70), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n581_), .B2(KEYINPUT12), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n499_), .A2(new_n579_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n485_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n560_), .A2(new_n592_), .A3(KEYINPUT12), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n496_), .A2(KEYINPUT68), .A3(new_n497_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT68), .B1(new_n496_), .B2(new_n497_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n579_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT70), .A3(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n590_), .A2(new_n591_), .A3(new_n593_), .A4(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n582_), .B(new_n588_), .C1(new_n599_), .C2(new_n578_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT69), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n513_), .A2(new_n519_), .A3(new_n505_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT65), .B1(new_n526_), .B2(new_n533_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n520_), .A2(new_n534_), .A3(KEYINPUT69), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n485_), .B1(new_n607_), .B2(new_n551_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n580_), .B1(new_n608_), .B2(KEYINPUT12), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n609_), .A2(new_n577_), .A3(new_n590_), .A4(new_n598_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n588_), .B1(new_n610_), .B2(new_n582_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n576_), .B1(new_n601_), .B2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n582_), .B1(new_n599_), .B2(new_n578_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n587_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(KEYINPUT72), .A3(new_n600_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n612_), .A2(KEYINPUT13), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT13), .B1(new_n612_), .B2(new_n615_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n456_), .A2(new_n457_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n538_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n458_), .A2(new_n557_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n458_), .B(new_n538_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT79), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT77), .B(G169gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT78), .B(G197gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n628_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n626_), .A2(new_n627_), .A3(new_n633_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n619_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n448_), .A2(new_n575_), .A3(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT101), .Z(new_n640_));
  INV_X1    g439(.A(new_n281_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n449_), .A3(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n643_));
  OR3_X1    g442(.A1(new_n642_), .A2(KEYINPUT103), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n643_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n448_), .A2(new_n638_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n571_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n504_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n281_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT103), .B1(new_n642_), .B2(new_n643_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n644_), .A2(new_n645_), .A3(new_n650_), .A4(new_n651_), .ZN(G1324gat));
  NOR3_X1   g451(.A1(new_n647_), .A2(new_n504_), .A3(new_n446_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n448_), .A2(new_n638_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n448_), .A2(KEYINPUT104), .A3(new_n638_), .A4(new_n653_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(G8gat), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n656_), .A2(KEYINPUT105), .A3(G8gat), .A4(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(KEYINPUT39), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(KEYINPUT39), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n662_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n660_), .A2(new_n663_), .A3(KEYINPUT39), .A4(new_n661_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n640_), .A2(new_n450_), .A3(new_n424_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .A4(new_n670_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1325gat));
  OR3_X1    g473(.A1(new_n639_), .A2(G15gat), .A3(new_n327_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n649_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n328_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(new_n677_), .B2(G15gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(G1326gat));
  OR3_X1    g480(.A1(new_n639_), .A2(G22gat), .A3(new_n444_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n676_), .A2(new_n381_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(G22gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n683_), .B2(G22gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n682_), .B1(new_n686_), .B2(new_n687_), .ZN(G1327gat));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n568_), .A2(new_n573_), .A3(new_n570_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n573_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n689_), .B1(new_n448_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n438_), .A2(new_n430_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n444_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n274_), .A2(KEYINPUT100), .A3(new_n276_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT100), .B1(new_n274_), .B2(new_n276_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n381_), .B(new_n446_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n328_), .B1(new_n695_), .B2(new_n698_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n281_), .A2(new_n328_), .A3(new_n425_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n689_), .B(new_n692_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n504_), .B(new_n638_), .C1(new_n693_), .C2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n699_), .A2(new_n700_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n572_), .A2(new_n574_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n701_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n705_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n710_), .A2(new_n504_), .A3(new_n638_), .A4(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(new_n641_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G29gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n504_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n571_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n448_), .A2(new_n638_), .A3(new_n716_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n281_), .A2(G29gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1328gat));
  NAND3_X1  g518(.A1(new_n706_), .A2(new_n424_), .A3(new_n712_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n717_), .A2(G36gat), .A3(new_n446_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT45), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(KEYINPUT45), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n721_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT46), .B1(new_n726_), .B2(KEYINPUT109), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n728_), .B(new_n729_), .C1(new_n721_), .C2(new_n725_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n727_), .A2(new_n730_), .ZN(G1329gat));
  NAND3_X1  g530(.A1(new_n706_), .A2(new_n328_), .A3(new_n712_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G43gat), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n717_), .A2(G43gat), .A3(new_n327_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(G1330gat));
  NAND3_X1  g536(.A1(new_n706_), .A2(new_n381_), .A3(new_n712_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G50gat), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n717_), .A2(G50gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n444_), .B2(new_n740_), .ZN(G1331gat));
  INV_X1    g540(.A(new_n637_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n618_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n707_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n648_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n746_), .A2(new_n461_), .A3(new_n281_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n575_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(KEYINPUT110), .A3(new_n575_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n641_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n461_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT111), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(new_n757_), .A3(new_n461_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n747_), .B1(new_n756_), .B2(new_n758_), .ZN(G1332gat));
  OAI21_X1  g558(.A(G64gat), .B1(new_n746_), .B2(new_n446_), .ZN(new_n760_));
  XOR2_X1   g559(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n424_), .A2(new_n462_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT113), .Z(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n752_), .B2(new_n764_), .ZN(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n746_), .B2(new_n327_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT49), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n328_), .A2(new_n470_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n752_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT114), .ZN(G1334gat));
  OAI21_X1  g569(.A(G78gat), .B1(new_n746_), .B2(new_n444_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT115), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT50), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n753_), .A2(new_n468_), .A3(new_n381_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1335gat));
  AOI211_X1 g574(.A(new_n715_), .B(new_n744_), .C1(new_n709_), .C2(new_n701_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n776_), .A2(new_n641_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n745_), .A2(new_n716_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n507_), .B1(new_n778_), .B2(new_n281_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1336gat));
  OAI21_X1  g579(.A(new_n384_), .B1(new_n778_), .B2(new_n446_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT116), .Z(new_n782_));
  NOR2_X1   g581(.A1(new_n446_), .A2(new_n384_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n776_), .B2(new_n783_), .ZN(G1337gat));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT117), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n527_), .B1(new_n776_), .B2(new_n328_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n778_), .A2(new_n518_), .A3(new_n327_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n785_), .A2(KEYINPUT117), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n789_), .B(new_n790_), .Z(G1338gat));
  NAND3_X1  g590(.A1(new_n710_), .A2(new_n504_), .A3(new_n743_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G106gat), .B1(new_n792_), .B2(new_n444_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n794_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n745_), .A2(new_n543_), .A3(new_n381_), .A4(new_n716_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT118), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n795_), .A2(new_n801_), .A3(new_n796_), .A4(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  NOR2_X1   g602(.A1(new_n626_), .A2(new_n634_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n621_), .A2(new_n623_), .ZN(new_n805_));
  MUX2_X1   g604(.A(new_n805_), .B(new_n625_), .S(new_n622_), .Z(new_n806_));
  AOI21_X1  g605(.A(new_n804_), .B1(new_n634_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n589_), .B(KEYINPUT12), .C1(new_n499_), .C2(new_n579_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT70), .B1(new_n596_), .B2(new_n597_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n577_), .B1(new_n812_), .B2(new_n609_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n610_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n599_), .A2(new_n814_), .A3(new_n578_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n588_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n637_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n814_), .B1(new_n599_), .B2(new_n578_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n599_), .A2(new_n578_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n587_), .B1(new_n823_), .B2(new_n816_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n819_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n601_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n809_), .B1(new_n820_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n647_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n612_), .A2(new_n615_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n807_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n600_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n587_), .B(new_n819_), .C1(new_n823_), .C2(new_n816_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n742_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n831_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT57), .B1(new_n835_), .B2(new_n571_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n829_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n601_), .B1(new_n818_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n808_), .B1(new_n824_), .B2(KEYINPUT56), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT58), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT120), .B1(new_n841_), .B2(new_n708_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n840_), .A3(KEYINPUT58), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n807_), .B1(new_n818_), .B2(new_n838_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n838_), .B(new_n587_), .C1(new_n823_), .C2(new_n816_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n600_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n692_), .A3(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n842_), .A2(new_n843_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n715_), .B1(new_n837_), .B2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n575_), .A2(new_n618_), .A3(new_n637_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n641_), .B(new_n328_), .C1(new_n852_), .C2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n425_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n742_), .ZN(new_n859_));
  INV_X1    g658(.A(G113gat), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n842_), .A2(new_n843_), .A3(new_n850_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n828_), .B1(new_n827_), .B2(new_n647_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n835_), .A2(KEYINPUT57), .A3(new_n571_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n504_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n853_), .B(KEYINPUT54), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n281_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n328_), .A4(new_n425_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT59), .B1(new_n856_), .B2(new_n857_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n870_), .A3(KEYINPUT121), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n860_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n859_), .B1(new_n875_), .B2(new_n742_), .ZN(G1340gat));
  OAI21_X1  g675(.A(G120gat), .B1(new_n871_), .B2(new_n618_), .ZN(new_n877_));
  INV_X1    g676(.A(G120gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n618_), .B2(KEYINPUT60), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n858_), .B(new_n879_), .C1(KEYINPUT60), .C2(new_n878_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n880_), .ZN(G1341gat));
  AOI21_X1  g680(.A(G127gat), .B1(new_n858_), .B2(new_n715_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(KEYINPUT122), .A2(G127gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G127gat), .B1(new_n504_), .B2(KEYINPUT122), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n882_), .B1(new_n884_), .B2(new_n885_), .ZN(G1342gat));
  AOI21_X1  g685(.A(G134gat), .B1(new_n858_), .B2(new_n647_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n873_), .A2(new_n874_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n692_), .A2(G134gat), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT123), .Z(new_n890_));
  AOI21_X1  g689(.A(new_n887_), .B1(new_n888_), .B2(new_n890_), .ZN(G1343gat));
  NAND4_X1  g690(.A1(new_n641_), .A2(new_n381_), .A3(new_n446_), .A4(new_n327_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(KEYINPUT124), .Z(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n742_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n619_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n715_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1346gat));
  AOI21_X1  g700(.A(G162gat), .B1(new_n894_), .B2(new_n647_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n894_), .A2(G162gat), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n904_), .B2(new_n692_), .ZN(G1347gat));
  XOR2_X1   g704(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n906_));
  NAND2_X1  g705(.A1(new_n865_), .A2(new_n866_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(new_n444_), .A3(new_n424_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n281_), .A3(new_n328_), .ZN(new_n910_));
  OAI211_X1 g709(.A(G169gat), .B(new_n906_), .C1(new_n910_), .C2(new_n637_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n906_), .ZN(new_n912_));
  NOR4_X1   g711(.A1(new_n908_), .A2(new_n641_), .A3(new_n637_), .A4(new_n327_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n301_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n304_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n911_), .A2(new_n914_), .A3(new_n915_), .ZN(G1348gat));
  NOR3_X1   g715(.A1(new_n908_), .A2(new_n641_), .A3(new_n327_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n619_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g718(.A1(new_n910_), .A2(new_n504_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n314_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(new_n290_), .B2(new_n920_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n910_), .B2(new_n708_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n917_), .A2(new_n647_), .A3(new_n395_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1351gat));
  NOR2_X1   g724(.A1(new_n446_), .A2(new_n328_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n907_), .A2(new_n445_), .A3(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n637_), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT126), .B(G197gat), .Z(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1352gat));
  INV_X1    g729(.A(new_n927_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n619_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n715_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  AND2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n934_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n937_), .B1(new_n934_), .B2(new_n935_), .ZN(G1354gat));
  NAND3_X1  g737(.A1(new_n931_), .A2(G218gat), .A3(new_n692_), .ZN(new_n939_));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n940_), .B1(new_n927_), .B2(new_n571_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n941_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


