//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n970_, new_n971_, new_n973_,
    new_n974_, new_n976_, new_n978_, new_n979_, new_n980_, new_n982_,
    new_n983_, new_n984_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT72), .B(G1gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n205_), .B1(new_n206_), .B2(G8gat), .ZN(new_n207_));
  INV_X1    g006(.A(G15gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(KEYINPUT71), .A2(G22gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT71), .A2(G22gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT71), .ZN(new_n212_));
  INV_X1    g011(.A(G22gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(KEYINPUT71), .A2(G22gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(G15gat), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT73), .B1(new_n207_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G1gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT72), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT72), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G1gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n222_), .A3(G8gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT14), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT73), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n216_), .A4(new_n211_), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n218_), .A2(new_n219_), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n219_), .B1(new_n218_), .B2(new_n226_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n204_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G1gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n218_), .A2(new_n219_), .A3(new_n226_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(G8gat), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G29gat), .A2(G36gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G29gat), .A2(G36gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(G43gat), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G29gat), .ZN(new_n238_));
  INV_X1    g037(.A(G36gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G43gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(new_n234_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n237_), .A2(new_n242_), .A3(G50gat), .ZN(new_n243_));
  AOI21_X1  g042(.A(G50gat), .B1(new_n237_), .B2(new_n242_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT76), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n229_), .A2(new_n233_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n203_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G169gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(G197gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(KEYINPUT77), .ZN(new_n254_));
  INV_X1    g053(.A(new_n246_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n227_), .A2(new_n228_), .A3(new_n204_), .ZN(new_n256_));
  AOI21_X1  g055(.A(G8gat), .B1(new_n231_), .B2(new_n232_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n244_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n237_), .A2(new_n242_), .A3(G50gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT15), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT15), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n229_), .A2(new_n233_), .A3(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n202_), .A3(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n249_), .A2(new_n254_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n254_), .B1(new_n249_), .B2(new_n266_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G57gat), .ZN(new_n270_));
  INV_X1    g069(.A(G64gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G57gat), .A2(G64gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G71gat), .B(G78gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT11), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n272_), .A2(new_n278_), .A3(new_n273_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n274_), .A2(new_n276_), .A3(KEYINPUT11), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G99gat), .A2(G106gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G85gat), .A2(G92gat), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT9), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G106gat), .ZN(new_n292_));
  INV_X1    g091(.A(G99gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT10), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT10), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G99gat), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n294_), .A2(new_n296_), .A3(KEYINPUT64), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT64), .B1(new_n294_), .B2(new_n296_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n292_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G85gat), .B(G92gat), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT9), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n291_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(new_n293_), .A3(new_n292_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n304_), .A2(new_n286_), .A3(new_n287_), .A4(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n300_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT8), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(KEYINPUT8), .A3(new_n300_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n283_), .B1(new_n302_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n291_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n313_), .A2(new_n309_), .A3(new_n310_), .A4(new_n282_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(KEYINPUT12), .A3(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n309_), .A2(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n313_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT12), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n283_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G230gat), .ZN(new_n321_));
  INV_X1    g120(.A(G233gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  OR3_X1    g124(.A1(new_n317_), .A2(KEYINPUT65), .A3(new_n283_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n312_), .A2(KEYINPUT65), .A3(new_n314_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G120gat), .B(G148gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G204gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT5), .ZN(new_n332_));
  INV_X1    g131(.A(G176gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n325_), .A2(new_n328_), .A3(new_n334_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(KEYINPUT13), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT13), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT66), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(KEYINPUT66), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n269_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n349_), .A2(new_n352_), .A3(new_n353_), .A4(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n360_), .A3(new_n357_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n362_), .A2(new_n350_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT85), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(G141gat), .B2(G148gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT85), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n361_), .A2(new_n363_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n359_), .A2(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(G127gat), .A2(G134gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G127gat), .A2(G134gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(G113gat), .A2(G120gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G113gat), .A2(G120gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n369_), .A2(new_n372_), .A3(new_n370_), .A4(new_n373_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT91), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT91), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n375_), .A2(new_n379_), .A3(new_n376_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n368_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n375_), .A2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n372_), .A2(new_n373_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n371_), .A2(new_n374_), .A3(KEYINPUT83), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n376_), .A2(KEYINPUT84), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n383_), .A2(new_n386_), .A3(new_n387_), .A4(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(new_n368_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT4), .B1(new_n381_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n389_), .A2(new_n368_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n391_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n368_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n392_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT0), .B(G57gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G85gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(G1gat), .B(G29gat), .Z(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n401_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT19), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n333_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G183gat), .A2(G190gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT23), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT79), .B(KEYINPUT23), .Z(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n415_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G183gat), .A2(G190gat), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n412_), .B(new_n414_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(KEYINPUT23), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n415_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n423_), .B(new_n424_), .C1(new_n417_), .C2(new_n415_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT25), .B(G183gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT26), .B(G190gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(G169gat), .A2(G176gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(KEYINPUT24), .A3(new_n412_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n429_), .A2(KEYINPUT24), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n425_), .A2(new_n428_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n420_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G197gat), .B(G204gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT21), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(G211gat), .A2(G218gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G211gat), .A2(G218gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G211gat), .B(G218gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT88), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n436_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n434_), .B(new_n435_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n442_), .A2(new_n440_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT20), .B1(new_n433_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n442_), .A2(new_n440_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n435_), .B2(new_n434_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n428_), .A2(new_n430_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT78), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT78), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n428_), .A2(new_n454_), .A3(new_n430_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n418_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .A4(new_n431_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n419_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n425_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n414_), .A2(KEYINPUT80), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n414_), .A2(KEYINPUT80), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n459_), .A2(new_n412_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n451_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n411_), .B1(new_n447_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT18), .B(G64gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G92gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G8gat), .B(G36gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n433_), .A2(new_n446_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT90), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n451_), .A3(new_n457_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n433_), .A2(new_n446_), .A3(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n470_), .A2(KEYINPUT20), .A3(new_n471_), .A4(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n464_), .B(new_n468_), .C1(new_n474_), .C2(new_n411_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(KEYINPUT20), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n478_), .A2(new_n410_), .A3(new_n470_), .A4(new_n473_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n468_), .B1(new_n479_), .B2(new_n464_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(KEYINPUT27), .ZN(new_n482_));
  INV_X1    g281(.A(new_n468_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n433_), .A2(new_n446_), .A3(new_n472_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n472_), .B1(new_n433_), .B2(new_n446_), .ZN(new_n485_));
  NOR4_X1   g284(.A1(new_n477_), .A2(new_n484_), .A3(new_n485_), .A4(new_n411_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n464_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n483_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n447_), .A2(new_n463_), .ZN(new_n489_));
  MUX2_X1   g288(.A(new_n489_), .B(new_n474_), .S(new_n411_), .Z(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n490_), .B2(new_n483_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT27), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n482_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT82), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n462_), .A2(new_n457_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT30), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n462_), .A2(new_n457_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n462_), .A2(new_n457_), .A3(new_n498_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n498_), .B1(new_n462_), .B2(new_n457_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n502_), .A2(new_n503_), .A3(KEYINPUT82), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G71gat), .B(G99gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G15gat), .B(G43gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n504_), .A2(KEYINPUT31), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT31), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n497_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n513_), .B2(new_n509_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n389_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n511_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT31), .B1(new_n504_), .B2(new_n510_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n512_), .A3(new_n509_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n389_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n501_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G78gat), .B(G106gat), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT29), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n359_), .B2(new_n367_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G228gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT86), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n446_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT86), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT87), .B1(new_n524_), .B2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n532_), .A2(new_n446_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n522_), .B(new_n530_), .C1(new_n533_), .C2(new_n526_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n368_), .A2(new_n523_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT28), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n368_), .A2(new_n539_), .A3(new_n523_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G22gat), .B(G50gat), .Z(new_n541_));
  AND3_X1   g340(.A1(new_n538_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n530_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n526_), .B1(new_n532_), .B2(new_n446_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n521_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n536_), .A2(new_n544_), .B1(new_n547_), .B2(new_n534_), .ZN(new_n548_));
  AND4_X1   g347(.A1(KEYINPUT89), .A2(new_n544_), .A3(new_n534_), .A4(new_n547_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n515_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n517_), .A2(new_n389_), .A3(new_n518_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n500_), .A3(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n520_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n550_), .B1(new_n520_), .B2(new_n553_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n408_), .B(new_n494_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT93), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n401_), .B2(new_n406_), .ZN(new_n559_));
  AOI211_X1 g358(.A(KEYINPUT33), .B(new_n405_), .C1(new_n397_), .C2(new_n400_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n488_), .B(new_n475_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n381_), .A2(new_n390_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n406_), .B1(new_n562_), .B2(new_n393_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT92), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n391_), .A2(new_n396_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n392_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(KEYINPUT92), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n564_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n557_), .B1(new_n561_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n483_), .A2(KEYINPUT32), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n571_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n407_), .B(new_n572_), .C1(new_n490_), .C2(new_n571_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n401_), .A2(new_n406_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT33), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n401_), .A2(new_n558_), .A3(new_n406_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n481_), .A2(new_n577_), .A3(KEYINPUT93), .A4(new_n568_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n570_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n520_), .A2(new_n553_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n550_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n556_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT70), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(G134gat), .ZN(new_n585_));
  INV_X1    g384(.A(G162gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n313_), .A2(new_n245_), .A3(new_n309_), .A4(new_n310_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT68), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT67), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT34), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT35), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n317_), .A2(new_n264_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n595_), .A2(KEYINPUT35), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n592_), .A2(new_n596_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n590_), .A2(new_n591_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n316_), .A2(new_n313_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n601_));
  OAI211_X1 g400(.A(KEYINPUT35), .B(new_n595_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n587_), .A2(new_n588_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n599_), .A2(new_n602_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n589_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n583_), .B1(new_n608_), .B2(KEYINPUT37), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n599_), .A2(new_n602_), .A3(new_n606_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n606_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n611_));
  OAI22_X1  g410(.A1(new_n610_), .A2(new_n611_), .B1(new_n588_), .B2(new_n587_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(KEYINPUT70), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT69), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(KEYINPUT69), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n609_), .A2(new_n614_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT16), .B(G183gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(G211gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT17), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n282_), .B(KEYINPUT74), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n229_), .A2(new_n233_), .A3(new_n625_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n628_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n229_), .A2(new_n233_), .A3(new_n625_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(new_n626_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT17), .B1(new_n630_), .B2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n624_), .B1(new_n634_), .B2(new_n622_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n630_), .A2(new_n633_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT75), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n638_), .B(new_n624_), .C1(new_n622_), .C2(new_n634_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n618_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n345_), .A2(new_n582_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n345_), .A2(new_n582_), .A3(KEYINPUT94), .A4(new_n643_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n206_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n407_), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT38), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n342_), .A2(new_n269_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n556_), .B2(new_n581_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n642_), .A2(new_n612_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n408_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n651_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n651_), .A2(KEYINPUT95), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1324gat));
  INV_X1    g461(.A(new_n494_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n646_), .A2(new_n204_), .A3(new_n663_), .A4(new_n647_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT96), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n665_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n654_), .A2(new_n655_), .A3(new_n663_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(new_n670_), .A3(G8gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G8gat), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n668_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT98), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT97), .B(KEYINPUT40), .Z(new_n677_));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n668_), .A2(new_n678_), .A3(new_n674_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n676_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n677_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n668_), .B2(new_n674_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT98), .B(new_n673_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n680_), .A2(new_n684_), .ZN(G1325gat));
  INV_X1    g484(.A(new_n580_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n648_), .A2(new_n208_), .A3(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT99), .Z(new_n688_));
  OAI21_X1  g487(.A(G15gat), .B1(new_n656_), .B2(new_n580_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT41), .Z(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1326gat));
  OAI21_X1  g490(.A(G22gat), .B1(new_n656_), .B2(new_n550_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT42), .ZN(new_n693_));
  INV_X1    g492(.A(new_n550_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n648_), .A2(new_n213_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1327gat));
  NAND2_X1  g495(.A1(new_n642_), .A2(new_n612_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT102), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n654_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n238_), .A3(new_n407_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT37), .B(new_n617_), .C1(new_n608_), .C2(KEYINPUT69), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n608_), .A2(new_n583_), .A3(KEYINPUT37), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT70), .B1(new_n612_), .B2(new_n613_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n556_), .B2(new_n581_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n642_), .B1(new_n706_), .B2(KEYINPUT43), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  AOI211_X1 g507(.A(new_n708_), .B(new_n705_), .C1(new_n556_), .C2(new_n581_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n707_), .A2(new_n653_), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT100), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n701_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n582_), .A2(new_n618_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n708_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n706_), .A2(KEYINPUT43), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n714_), .A2(new_n642_), .A3(new_n652_), .A4(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(KEYINPUT100), .A3(KEYINPUT44), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n712_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n238_), .B1(new_n718_), .B2(new_n407_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT101), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT101), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n700_), .B1(new_n720_), .B2(new_n721_), .ZN(G1328gat));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n239_), .B1(new_n718_), .B2(new_n663_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n699_), .A2(new_n239_), .A3(new_n663_), .ZN(new_n725_));
  XOR2_X1   g524(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n723_), .B(KEYINPUT46), .C1(new_n724_), .C2(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n710_), .A2(new_n711_), .A3(new_n701_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT44), .B1(new_n716_), .B2(KEYINPUT100), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n663_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G36gat), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n723_), .A2(KEYINPUT46), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n723_), .A2(KEYINPUT46), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .A4(new_n727_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n729_), .A2(new_n736_), .ZN(G1329gat));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n718_), .A2(new_n686_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G43gat), .ZN(new_n740_));
  INV_X1    g539(.A(new_n699_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n741_), .A2(G43gat), .A3(new_n580_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n738_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT47), .B(new_n742_), .C1(new_n739_), .C2(G43gat), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1330gat));
  NAND3_X1  g545(.A1(new_n718_), .A2(G50gat), .A3(new_n694_), .ZN(new_n747_));
  INV_X1    g546(.A(G50gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n741_), .B2(new_n550_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(G1331gat));
  INV_X1    g551(.A(new_n269_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n556_), .B2(new_n581_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n343_), .A2(new_n344_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n655_), .A3(new_n755_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n756_), .A2(new_n270_), .A3(new_n408_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n754_), .B(KEYINPUT106), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n342_), .A3(new_n643_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n759_), .A2(new_n408_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(new_n760_), .B2(new_n270_), .ZN(G1332gat));
  OAI21_X1  g560(.A(G64gat), .B1(new_n756_), .B2(new_n494_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT48), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n663_), .A2(new_n271_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n759_), .B2(new_n764_), .ZN(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n756_), .B2(new_n580_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT49), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n759_), .A2(G71gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n580_), .ZN(G1334gat));
  OAI21_X1  g568(.A(G78gat), .B1(new_n756_), .B2(new_n550_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT50), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n759_), .A2(G78gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n550_), .ZN(G1335gat));
  NAND3_X1  g572(.A1(new_n758_), .A2(new_n755_), .A3(new_n698_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(new_n408_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n707_), .A2(new_n709_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n342_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(new_n753_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n407_), .ZN(new_n780_));
  MUX2_X1   g579(.A(new_n775_), .B(new_n780_), .S(G85gat), .Z(G1336gat));
  INV_X1    g580(.A(G92gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n774_), .B2(new_n494_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT107), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n494_), .A2(new_n782_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n779_), .B2(new_n785_), .ZN(G1337gat));
  NOR2_X1   g585(.A1(new_n297_), .A2(new_n298_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n774_), .A2(new_n787_), .A3(new_n580_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n293_), .B1(new_n779_), .B2(new_n686_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT51), .Z(G1338gat));
  OR3_X1    g590(.A1(new_n774_), .A2(G106gat), .A3(new_n550_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n776_), .A2(new_n694_), .A3(new_n778_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G106gat), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n793_), .A3(G106gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT53), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n792_), .B(new_n799_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1339gat));
  NAND2_X1  g600(.A1(new_n494_), .A2(new_n407_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n554_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(KEYINPUT112), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(KEYINPUT112), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT59), .ZN(new_n807_));
  INV_X1    g606(.A(new_n642_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n337_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT108), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT111), .B1(new_n812_), .B2(KEYINPUT110), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT55), .B1(new_n320_), .B2(new_n324_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n323_), .A2(KEYINPUT109), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n320_), .B2(KEYINPUT55), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  INV_X1    g616(.A(new_n815_), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n817_), .B(new_n818_), .C1(new_n315_), .C2(new_n319_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n814_), .A2(new_n816_), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n813_), .B1(new_n820_), .B2(new_n334_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n337_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n325_), .A2(new_n817_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n320_), .A2(KEYINPUT55), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n818_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n320_), .A2(KEYINPUT55), .A3(new_n815_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n813_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n812_), .A2(KEYINPUT111), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n828_), .A2(new_n335_), .A3(new_n829_), .A4(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n811_), .A2(new_n821_), .A3(new_n823_), .A4(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n258_), .A2(new_n265_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n203_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n229_), .A2(new_n233_), .A3(new_n246_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n258_), .A2(new_n202_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n253_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n249_), .A2(new_n253_), .A3(new_n266_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n338_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n809_), .B(new_n612_), .C1(new_n832_), .C2(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n820_), .A2(new_n812_), .A3(new_n334_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n335_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n337_), .B(new_n839_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n812_), .B1(new_n820_), .B2(new_n334_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n335_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n849_), .A2(KEYINPUT58), .A3(new_n337_), .A4(new_n839_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n846_), .A2(new_n618_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n612_), .B1(new_n832_), .B2(new_n840_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(KEYINPUT57), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n841_), .B1(new_n853_), .B2(KEYINPUT113), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n851_), .B(new_n855_), .C1(new_n852_), .C2(KEYINPUT57), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n808_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n643_), .A2(new_n858_), .A3(new_n269_), .A4(new_n777_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n705_), .A2(new_n640_), .A3(new_n641_), .A4(new_n269_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT54), .B1(new_n860_), .B2(new_n342_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n807_), .B1(new_n857_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT114), .ZN(new_n864_));
  INV_X1    g663(.A(G113gat), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n269_), .A2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n642_), .B1(new_n853_), .B2(new_n841_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n859_), .A2(new_n861_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n804_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT59), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n807_), .B(new_n872_), .C1(new_n857_), .C2(new_n862_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n864_), .A2(new_n866_), .A3(new_n871_), .A4(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n865_), .B1(new_n870_), .B2(new_n269_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT115), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n874_), .A2(new_n878_), .A3(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1340gat));
  INV_X1    g679(.A(new_n870_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT116), .B(G120gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n777_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(KEYINPUT60), .B2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(KEYINPUT60), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n882_), .ZN(new_n886_));
  AND4_X1   g685(.A1(new_n871_), .A2(new_n884_), .A3(new_n864_), .A4(new_n873_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n755_), .ZN(G1341gat));
  AOI21_X1  g687(.A(G127gat), .B1(new_n881_), .B2(new_n808_), .ZN(new_n889_));
  AND4_X1   g688(.A1(G127gat), .A2(new_n864_), .A3(new_n871_), .A4(new_n873_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n808_), .ZN(G1342gat));
  AOI21_X1  g690(.A(G134gat), .B1(new_n881_), .B2(new_n612_), .ZN(new_n892_));
  AND4_X1   g691(.A1(G134gat), .A2(new_n864_), .A3(new_n871_), .A4(new_n873_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n618_), .ZN(G1343gat));
  AND2_X1   g693(.A1(new_n869_), .A2(new_n555_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n802_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n269_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n347_), .ZN(G1344gat));
  AND2_X1   g698(.A1(new_n895_), .A2(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n755_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT117), .B(G148gat), .Z(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1345gat));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n900_), .A2(new_n808_), .A3(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n897_), .B2(new_n642_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n906_), .A2(new_n909_), .A3(new_n907_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1346gat));
  OAI21_X1  g712(.A(new_n586_), .B1(new_n897_), .B2(new_n608_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n618_), .A2(G162gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n897_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n914_), .B(KEYINPUT120), .C1(new_n897_), .C2(new_n915_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n494_), .A2(new_n407_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n803_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n753_), .B(new_n923_), .C1(new_n857_), .C2(new_n862_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G169gat), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n924_), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n927_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n923_), .B1(new_n857_), .B2(new_n862_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT123), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n933_), .B(new_n923_), .C1(new_n857_), .C2(new_n862_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n753_), .A2(new_n413_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT124), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n930_), .B(new_n938_), .C1(new_n927_), .C2(new_n929_), .ZN(G1348gat));
  AOI21_X1  g738(.A(new_n694_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n922_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n832_), .A2(new_n840_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n608_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n809_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n852_), .A2(KEYINPUT57), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n945_), .A2(new_n946_), .A3(new_n851_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n862_), .B1(new_n947_), .B2(new_n642_), .ZN(new_n948_));
  OAI21_X1  g747(.A(KEYINPUT125), .B1(new_n948_), .B2(new_n694_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n942_), .A2(new_n949_), .A3(new_n686_), .A4(new_n755_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n950_), .A2(G176gat), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n342_), .A2(new_n333_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n952_), .B1(new_n932_), .B2(new_n934_), .ZN(new_n953_));
  OAI21_X1  g752(.A(KEYINPUT126), .B1(new_n951_), .B2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n950_), .A2(G176gat), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956_));
  AND2_X1   g755(.A1(new_n932_), .A2(new_n934_), .ZN(new_n957_));
  OAI211_X1 g756(.A(new_n955_), .B(new_n956_), .C1(new_n957_), .C2(new_n952_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n954_), .A2(new_n958_), .ZN(G1349gat));
  NAND4_X1  g758(.A1(new_n942_), .A2(new_n949_), .A3(new_n808_), .A4(new_n686_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(new_n962_));
  AOI211_X1 g761(.A(new_n580_), .B(new_n922_), .C1(new_n940_), .C2(new_n941_), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n963_), .A2(KEYINPUT127), .A3(new_n808_), .A4(new_n949_), .ZN(new_n964_));
  INV_X1    g763(.A(G183gat), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n962_), .A2(new_n964_), .A3(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n426_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n935_), .A2(new_n808_), .A3(new_n967_), .ZN(new_n968_));
  AND2_X1   g767(.A1(new_n966_), .A2(new_n968_), .ZN(G1350gat));
  OAI21_X1  g768(.A(G190gat), .B1(new_n957_), .B2(new_n705_), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n935_), .A2(new_n612_), .A3(new_n427_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(G1351gat));
  AND2_X1   g771(.A1(new_n895_), .A2(new_n921_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(new_n753_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g774(.A1(new_n973_), .A2(new_n755_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g776(.A1(new_n973_), .A2(new_n808_), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n978_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n979_));
  XOR2_X1   g778(.A(KEYINPUT63), .B(G211gat), .Z(new_n980_));
  OAI21_X1  g779(.A(new_n979_), .B1(new_n978_), .B2(new_n980_), .ZN(G1354gat));
  AOI21_X1  g780(.A(G218gat), .B1(new_n973_), .B2(new_n612_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n618_), .A2(G218gat), .ZN(new_n983_));
  INV_X1    g782(.A(new_n983_), .ZN(new_n984_));
  AOI21_X1  g783(.A(new_n982_), .B1(new_n973_), .B2(new_n984_), .ZN(G1355gat));
endmodule


