//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_;
  XNOR2_X1  g000(.A(G1gat), .B(G8gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G15gat), .A2(G22gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G1gat), .A2(G8gat), .ZN(new_n207_));
  AOI22_X1  g006(.A1(new_n205_), .A2(new_n206_), .B1(KEYINPUT14), .B2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n204_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(G43gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(G43gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(G50gat), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(G50gat), .B1(new_n211_), .B2(new_n212_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT81), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n209_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(new_n209_), .B2(new_n216_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n216_), .A2(KEYINPUT15), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n209_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n221_), .A2(new_n231_), .A3(new_n223_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G141gat), .ZN(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G197gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n225_), .A2(new_n232_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n225_), .B2(new_n232_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G120gat), .B(G148gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G176gat), .B(G204gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G230gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT8), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G99gat), .A2(G106gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT6), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(G99gat), .ZN(new_n259_));
  INV_X1    g058(.A(G106gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT7), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G99gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(new_n260_), .A3(KEYINPUT64), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT7), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n257_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n252_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n256_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT7), .B1(new_n259_), .B2(new_n260_), .ZN(new_n272_));
  AND4_X1   g071(.A1(KEYINPUT64), .A2(new_n262_), .A3(new_n260_), .A4(KEYINPUT7), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n271_), .B(new_n267_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(G85gat), .A2(G92gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G85gat), .A2(G92gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT66), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G85gat), .ZN(new_n278_));
  INV_X1    g077(.A(G92gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G85gat), .A2(G92gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n274_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT67), .B1(new_n268_), .B2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n277_), .A2(new_n283_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n267_), .B2(new_n266_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT8), .B1(new_n289_), .B2(KEYINPUT65), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT68), .B1(new_n266_), .B2(new_n287_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n294_), .A3(new_n284_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(KEYINPUT8), .A3(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n286_), .A2(new_n292_), .A3(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n275_), .A2(new_n276_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n257_), .B1(new_n298_), .B2(KEYINPUT9), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT10), .B(G99gat), .ZN(new_n300_));
  OAI221_X1 g099(.A(new_n299_), .B1(KEYINPUT9), .B2(new_n282_), .C1(G106gat), .C2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G57gat), .B(G64gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT69), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G71gat), .B(G78gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(KEYINPUT11), .A3(new_n307_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n297_), .A3(new_n301_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(KEYINPUT12), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT12), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n302_), .A2(new_n312_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n251_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n250_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n249_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n317_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n250_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n319_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n248_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n318_), .A2(new_n319_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT71), .B1(new_n327_), .B2(new_n248_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n320_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT13), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n325_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(KEYINPUT71), .A3(new_n248_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT13), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n320_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G127gat), .B(G155gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G183gat), .B(G211gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT17), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G231gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n311_), .B(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n345_), .A2(new_n230_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n230_), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT17), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n343_), .B1(new_n348_), .B2(new_n341_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n347_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT79), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n351_), .B(new_n343_), .C1(new_n341_), .C2(new_n348_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT74), .B(G190gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G218gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G134gat), .B(G162gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT36), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G232gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT72), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT34), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT35), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n297_), .A2(new_n216_), .A3(new_n301_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n297_), .A2(KEYINPUT73), .A3(new_n216_), .A4(new_n301_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n364_), .A2(new_n365_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n297_), .A2(new_n301_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AND4_X1   g174(.A1(new_n367_), .A2(new_n372_), .A3(new_n373_), .A4(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n367_), .B1(new_n377_), .B2(new_n373_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n360_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n366_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n367_), .A3(new_n373_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT36), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n359_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT75), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(KEYINPUT76), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(KEYINPUT37), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT37), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n379_), .B(new_n386_), .C1(KEYINPUT76), .C2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n355_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n336_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT80), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT97), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G204gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G197gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n236_), .A2(G204gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT90), .ZN(new_n402_));
  OR3_X1    g201(.A1(new_n236_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(KEYINPUT21), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G211gat), .B(G218gat), .Z(new_n407_));
  INV_X1    g206(.A(KEYINPUT21), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n400_), .A2(new_n401_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n402_), .A2(new_n403_), .A3(KEYINPUT91), .A4(KEYINPUT21), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT25), .B(G183gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT26), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G190gat), .ZN(new_n415_));
  INV_X1    g214(.A(G190gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT26), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n415_), .A2(new_n417_), .A3(KEYINPUT95), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT95), .B1(new_n415_), .B2(new_n417_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n413_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT23), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(G183gat), .B2(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(KEYINPUT23), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n421_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n421_), .B1(new_n424_), .B2(KEYINPUT23), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G176gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT24), .B1(new_n234_), .B2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432_));
  MUX2_X1   g231(.A(new_n431_), .B(KEYINPUT24), .S(new_n432_), .Z(new_n433_));
  NAND3_X1  g232(.A1(new_n420_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n408_), .B1(new_n407_), .B2(KEYINPUT92), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G211gat), .B(G218gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT92), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n409_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n424_), .B(KEYINPUT23), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(G183gat), .B2(G190gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n234_), .A2(new_n430_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT22), .B(G169gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(new_n430_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n412_), .A2(new_n434_), .A3(new_n440_), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT20), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n427_), .B1(new_n441_), .B2(new_n421_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT82), .B(G190gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(G183gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n445_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n415_), .B(new_n413_), .C1(new_n450_), .C2(new_n414_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n433_), .A2(new_n441_), .A3(new_n453_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n452_), .A2(new_n454_), .B1(new_n412_), .B2(new_n440_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n398_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G64gat), .B(G92gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n412_), .A2(new_n440_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n434_), .A2(new_n446_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n452_), .A2(new_n412_), .A3(new_n440_), .A4(new_n454_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n464_), .A2(KEYINPUT20), .A3(new_n465_), .A4(new_n397_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n456_), .A2(new_n461_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n461_), .B1(new_n456_), .B2(new_n466_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n395_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n456_), .A2(new_n466_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n461_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n456_), .A2(new_n461_), .A3(new_n466_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(KEYINPUT97), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G141gat), .A2(G148gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n476_), .B(KEYINPUT86), .Z(new_n477_));
  NAND2_X1  g276(.A1(G141gat), .A2(G148gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(G155gat), .B(G162gat), .Z(new_n479_));
  INV_X1    g278(.A(KEYINPUT1), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n477_), .A2(new_n478_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT2), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT2), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n478_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT3), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n476_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n486_), .A2(new_n488_), .A3(new_n489_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n479_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n492_), .B2(new_n479_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n483_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(G127gat), .A2(G134gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G127gat), .A2(G134gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G113gat), .ZN(new_n500_));
  INV_X1    g299(.A(G113gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n501_), .A3(new_n498_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n500_), .A2(G120gat), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(G120gat), .B1(new_n500_), .B2(new_n502_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n496_), .A2(new_n506_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n505_), .B(new_n483_), .C1(new_n495_), .C2(new_n494_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G225gat), .A2(G233gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(KEYINPUT4), .A3(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n510_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT4), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n496_), .A2(new_n506_), .A3(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT0), .B(G57gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(G85gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(G1gat), .B(G29gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n511_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n511_), .A2(new_n516_), .A3(new_n520_), .A4(new_n522_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n509_), .A2(new_n513_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n512_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n520_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n475_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT99), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n471_), .A2(KEYINPUT32), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n470_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n511_), .A2(new_n516_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n529_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n397_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n464_), .A2(KEYINPUT20), .A3(new_n465_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(new_n397_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n533_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n536_), .A2(new_n521_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n492_), .A2(new_n479_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT88), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n492_), .A2(new_n493_), .A3(new_n479_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n481_), .A2(new_n478_), .A3(new_n482_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n543_), .A2(new_n544_), .B1(new_n545_), .B2(new_n477_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G22gat), .B(G50gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT28), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n496_), .B2(KEYINPUT29), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n462_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G228gat), .A2(G233gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT89), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n462_), .B(new_n556_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n553_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G78gat), .B(G106gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(KEYINPUT94), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n561_), .B(KEYINPUT93), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n563_), .A2(new_n565_), .A3(new_n559_), .A4(new_n558_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n553_), .A2(KEYINPUT94), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n558_), .A2(new_n565_), .A3(new_n559_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n565_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n534_), .A2(new_n541_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT99), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n475_), .A2(new_n526_), .A3(new_n574_), .A4(new_n530_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n532_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n452_), .A2(new_n454_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT30), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT85), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n452_), .A2(new_n580_), .A3(new_n454_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G71gat), .B(G99gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(G43gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT84), .B(G15gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G227gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n585_), .B(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n582_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n583_), .B1(new_n582_), .B2(new_n589_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n505_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n582_), .A2(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT31), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n506_), .A3(new_n590_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n579_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n593_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n539_), .A2(new_n461_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(KEYINPUT27), .A3(new_n472_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT100), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n536_), .A2(new_n521_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT27), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n603_), .A2(new_n609_), .A3(new_n472_), .A4(KEYINPUT27), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n605_), .A2(new_n606_), .A3(new_n608_), .A4(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n562_), .B(new_n566_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n602_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n576_), .A2(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n593_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n598_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n606_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n605_), .A2(new_n612_), .A3(new_n608_), .A4(new_n610_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT80), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n336_), .A2(new_n392_), .A3(new_n623_), .ZN(new_n624_));
  AND4_X1   g423(.A1(new_n243_), .A2(new_n394_), .A3(new_n622_), .A4(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(G1gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n606_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n336_), .A2(new_n243_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n620_), .B1(new_n576_), .B2(new_n614_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n387_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n355_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n637_), .B2(new_n606_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n628_), .A2(new_n629_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n630_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(G1324gat));
  AND2_X1   g441(.A1(new_n605_), .A2(new_n610_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(new_n608_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n636_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G8gat), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(KEYINPUT39), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(KEYINPUT39), .ZN(new_n649_));
  INV_X1    g448(.A(new_n625_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n644_), .A2(G8gat), .ZN(new_n651_));
  OAI22_X1  g450(.A1(new_n648_), .A2(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(G1325gat));
  INV_X1    g453(.A(new_n602_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G15gat), .B1(new_n637_), .B2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT41), .Z(new_n657_));
  OR2_X1    g456(.A1(new_n655_), .A2(G15gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n650_), .B2(new_n658_), .ZN(G1326gat));
  OAI21_X1  g458(.A(G22gat), .B1(new_n637_), .B2(new_n612_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n612_), .A2(G22gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT102), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n650_), .B2(new_n663_), .ZN(G1327gat));
  AOI21_X1  g463(.A(new_n242_), .B1(new_n330_), .B2(new_n335_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n389_), .A2(KEYINPUT104), .A3(new_n391_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT104), .B1(new_n389_), .B2(new_n391_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n666_), .B1(new_n669_), .B2(new_n622_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n389_), .A2(new_n391_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n632_), .A2(KEYINPUT43), .A3(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n355_), .B(new_n665_), .C1(new_n670_), .C2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G29gat), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n671_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n389_), .A2(KEYINPUT104), .A3(new_n391_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n622_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n666_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n672_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n684_), .A2(KEYINPUT44), .A3(new_n355_), .A4(new_n665_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n627_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n355_), .A2(new_n634_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT105), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(new_n665_), .A3(new_n622_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n606_), .ZN(new_n691_));
  OAI22_X1  g490(.A1(new_n676_), .A2(new_n686_), .B1(G29gat), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT106), .ZN(G1328gat));
  XNOR2_X1  g492(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695_));
  INV_X1    g494(.A(G36gat), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n689_), .A2(new_n695_), .A3(new_n696_), .A4(new_n645_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n633_), .A2(new_n696_), .A3(new_n688_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT107), .B1(new_n698_), .B2(new_n644_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n699_), .A3(KEYINPUT45), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n675_), .A2(new_n645_), .A3(new_n685_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n694_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n707_));
  AND4_X1   g506(.A1(new_n694_), .A2(new_n706_), .A3(new_n703_), .A4(new_n702_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710_));
  AOI21_X1  g509(.A(G43gat), .B1(new_n689_), .B2(new_n602_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n672_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n355_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n631_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n655_), .B1(new_n714_), .B2(KEYINPUT44), .ZN(new_n715_));
  INV_X1    g514(.A(G43gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT109), .B(new_n711_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n675_), .A2(G43gat), .A3(new_n602_), .A4(new_n685_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n711_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n710_), .B1(new_n718_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G43gat), .B1(new_n714_), .B2(KEYINPUT44), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n685_), .A2(new_n602_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT109), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n720_), .A2(new_n719_), .A3(new_n721_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(KEYINPUT47), .A3(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n723_), .A2(new_n729_), .ZN(G1330gat));
  NAND3_X1  g529(.A1(new_n675_), .A2(new_n613_), .A3(new_n685_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G50gat), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n612_), .A2(G50gat), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT110), .Z(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n690_), .B2(new_n734_), .ZN(G1331gat));
  NOR2_X1   g534(.A1(new_n336_), .A2(new_n243_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n622_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n635_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(G57gat), .A3(new_n627_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT111), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(KEYINPUT111), .ZN(new_n743_));
  INV_X1    g542(.A(new_n671_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n737_), .A2(new_n355_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G57gat), .B1(new_n745_), .B2(new_n627_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n742_), .A2(new_n743_), .A3(new_n746_), .ZN(G1332gat));
  NAND3_X1  g546(.A1(new_n738_), .A2(new_n635_), .A3(new_n645_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(G64gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G64gat), .ZN(new_n751_));
  INV_X1    g550(.A(new_n745_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n644_), .A2(G64gat), .ZN(new_n753_));
  OAI22_X1  g552(.A1(new_n750_), .A2(new_n751_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT112), .ZN(G1333gat));
  OR3_X1    g554(.A1(new_n752_), .A2(G71gat), .A3(new_n655_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n740_), .A2(new_n602_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(G71gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G71gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n740_), .A2(new_n613_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G78gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G78gat), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n766_));
  OR3_X1    g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n612_), .A2(G78gat), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT114), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n767_), .B(new_n768_), .C1(new_n752_), .C2(new_n770_), .ZN(G1335gat));
  AND2_X1   g570(.A1(new_n738_), .A2(new_n688_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n627_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n684_), .A2(new_n355_), .A3(new_n736_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n627_), .A2(G85gat), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT115), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n773_), .B1(new_n775_), .B2(new_n777_), .ZN(G1336gat));
  NOR3_X1   g577(.A1(new_n774_), .A2(new_n279_), .A3(new_n644_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G92gat), .B1(new_n772_), .B2(new_n645_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n774_), .B2(new_n655_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n300_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n772_), .A2(new_n783_), .A3(new_n602_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n772_), .A2(new_n260_), .A3(new_n613_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G106gat), .B1(new_n774_), .B2(new_n612_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(KEYINPUT52), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(KEYINPUT52), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n787_), .B(new_n793_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  NAND3_X1  g594(.A1(new_n336_), .A2(new_n392_), .A3(new_n242_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n336_), .A2(new_n392_), .A3(KEYINPUT54), .A4(new_n242_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT116), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n321_), .A2(new_n250_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n322_), .A2(KEYINPUT55), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n318_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n803_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n802_), .B1(new_n807_), .B2(new_n248_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n318_), .A2(new_n805_), .ZN(new_n809_));
  AOI211_X1 g608(.A(KEYINPUT55), .B(new_n251_), .C1(new_n315_), .C2(new_n317_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n809_), .A2(new_n810_), .B1(new_n250_), .B2(new_n321_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n811_), .A2(KEYINPUT116), .A3(new_n801_), .A4(new_n249_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n242_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n808_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n221_), .A2(new_n231_), .A3(KEYINPUT117), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT117), .B1(new_n221_), .B2(new_n231_), .ZN(new_n817_));
  OR3_X1    g616(.A1(new_n816_), .A2(new_n223_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n222_), .A2(new_n223_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n237_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n239_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n329_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n814_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n387_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n811_), .A2(new_n249_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n811_), .A2(new_n801_), .A3(new_n249_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n829_), .A2(new_n333_), .A3(new_n822_), .A4(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n821_), .B1(new_n828_), .B2(KEYINPUT56), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(KEYINPUT58), .A3(new_n333_), .A4(new_n830_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n835_), .A3(new_n744_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n824_), .A2(KEYINPUT57), .A3(new_n387_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n827_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n800_), .B1(new_n838_), .B2(new_n355_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n644_), .A2(new_n627_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n840_), .A2(new_n613_), .A3(new_n655_), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n841_), .B(KEYINPUT118), .Z(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT119), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n634_), .B1(new_n814_), .B2(new_n823_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(new_n826_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n713_), .B1(new_n847_), .B2(new_n836_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n845_), .B(new_n842_), .C1(new_n848_), .C2(new_n800_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n844_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850_), .B2(new_n243_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(KEYINPUT120), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(KEYINPUT120), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n838_), .A2(new_n355_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n800_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n860_), .B2(new_n842_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n839_), .A2(new_n843_), .A3(new_n855_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n852_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n856_), .B(new_n855_), .C1(new_n839_), .C2(new_n843_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(new_n842_), .A3(new_n854_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(KEYINPUT121), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n242_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n851_), .B1(new_n867_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g667(.A(new_n336_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G120gat), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n872_));
  AOI21_X1  g671(.A(G120gat), .B1(new_n869_), .B2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n844_), .B2(new_n849_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(G120gat), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n874_), .A2(KEYINPUT122), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT122), .B1(new_n874_), .B2(new_n875_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n871_), .B1(new_n876_), .B2(new_n877_), .ZN(G1341gat));
  AOI21_X1  g677(.A(G127gat), .B1(new_n850_), .B2(new_n713_), .ZN(new_n879_));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n881_), .B2(new_n713_), .ZN(G1342gat));
  AOI21_X1  g681(.A(G134gat), .B1(new_n850_), .B2(new_n634_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT123), .B(G134gat), .Z(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n885_), .B2(new_n744_), .ZN(G1343gat));
  NOR2_X1   g685(.A1(new_n602_), .A2(new_n612_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n839_), .A2(new_n840_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n243_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT124), .B(G141gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1344gat));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n869_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n713_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  AOI21_X1  g696(.A(G162gat), .B1(new_n889_), .B2(new_n634_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n669_), .A2(G162gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n889_), .B2(new_n899_), .ZN(G1347gat));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n839_), .A2(new_n613_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n644_), .A2(new_n627_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n602_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n242_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n901_), .B1(new_n907_), .B2(new_n234_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n444_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT62), .B(G169gat), .C1(new_n906_), .C2(new_n242_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .ZN(G1348gat));
  INV_X1    g710(.A(new_n906_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G176gat), .B1(new_n912_), .B2(new_n869_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n860_), .A2(new_n612_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n904_), .B1(new_n914_), .B2(KEYINPUT125), .ZN(new_n915_));
  OR3_X1    g714(.A1(new_n839_), .A2(KEYINPUT125), .A3(new_n613_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n915_), .A2(G176gat), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n913_), .B1(new_n917_), .B2(new_n869_), .ZN(G1349gat));
  NOR3_X1   g717(.A1(new_n906_), .A2(new_n355_), .A3(new_n413_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n915_), .A2(new_n713_), .A3(new_n916_), .ZN(new_n920_));
  INV_X1    g719(.A(G183gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(G1350gat));
  OR2_X1    g721(.A1(new_n418_), .A2(new_n419_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n902_), .A2(new_n634_), .A3(new_n923_), .A4(new_n905_), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n839_), .A2(new_n613_), .A3(new_n671_), .A4(new_n904_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n416_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n924_), .B(KEYINPUT126), .C1(new_n416_), .C2(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1351gat));
  NAND3_X1  g729(.A1(new_n860_), .A2(new_n887_), .A3(new_n903_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n242_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n236_), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n336_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(new_n399_), .ZN(G1353gat));
  AOI21_X1  g734(.A(new_n355_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT127), .B1(new_n931_), .B2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n839_), .A2(new_n888_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n940_), .A2(new_n941_), .A3(new_n903_), .A4(new_n936_), .ZN(new_n942_));
  AND3_X1   g741(.A1(new_n938_), .A2(new_n939_), .A3(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n939_), .B1(new_n938_), .B2(new_n942_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1354gat));
  INV_X1    g744(.A(G218gat), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n931_), .A2(new_n946_), .A3(new_n671_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n940_), .A2(new_n634_), .A3(new_n903_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n946_), .ZN(G1355gat));
endmodule


