//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n205_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(G231gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT77), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  INV_X1    g012(.A(G8gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G1gat), .B(G8gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n212_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G127gat), .B(G155gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT16), .ZN(new_n222_));
  XOR2_X1   g021(.A(G183gat), .B(G211gat), .Z(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n219_), .B1(new_n220_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(KEYINPUT17), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(new_n219_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT78), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G29gat), .B(G36gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n230_), .A2(KEYINPUT70), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(KEYINPUT70), .ZN(new_n232_));
  XOR2_X1   g031(.A(G43gat), .B(G50gat), .Z(new_n233_));
  OR3_X1    g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(new_n218_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n236_), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n218_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n236_), .A2(new_n218_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n238_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n240_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G113gat), .B(G141gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G169gat), .B(G197gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n251_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G99gat), .A2(G106gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT6), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT6), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(G99gat), .A3(G106gat), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G106gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT10), .B(G99gat), .Z(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G85gat), .ZN(new_n265_));
  INV_X1    g064(.A(G92gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT9), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G85gat), .A2(G92gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n268_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n269_), .B2(new_n268_), .ZN(new_n272_));
  OAI221_X1 g071(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n264_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT8), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT7), .ZN(new_n276_));
  INV_X1    g075(.A(G99gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n262_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT65), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n258_), .A2(new_n260_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(new_n283_), .A3(new_n279_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n267_), .A2(new_n269_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n275_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n275_), .B(new_n287_), .C1(new_n261_), .C2(new_n280_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n274_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(KEYINPUT66), .B(new_n274_), .C1(new_n288_), .C2(new_n290_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n209_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n209_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G230gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT67), .B1(new_n288_), .B2(new_n290_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n280_), .A2(KEYINPUT65), .B1(new_n258_), .B2(new_n260_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n286_), .B1(new_n307_), .B2(new_n284_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n306_), .B(new_n289_), .C1(new_n308_), .C2(new_n275_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n274_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n297_), .A2(KEYINPUT12), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n304_), .A2(new_n314_), .A3(new_n296_), .A4(new_n300_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT5), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G176gat), .B(G204gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n302_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(new_n302_), .B2(new_n315_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT13), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n324_), .B1(KEYINPUT69), .B2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n229_), .A2(new_n256_), .A3(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT100), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337_));
  INV_X1    g136(.A(G141gat), .ZN(new_n338_));
  INV_X1    g137(.A(G148gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT84), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(KEYINPUT84), .A3(new_n337_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n336_), .B1(new_n345_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n346_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n334_), .B1(KEYINPUT1), .B2(new_n332_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n332_), .A2(KEYINPUT1), .ZN(new_n356_));
  AOI211_X1 g155(.A(new_n343_), .B(new_n354_), .C1(new_n355_), .C2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT29), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G197gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G204gat), .ZN(new_n360_));
  INV_X1    g159(.A(G204gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G197gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT21), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G211gat), .B(G218gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n361_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n359_), .A2(G204gat), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT21), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT85), .B1(new_n361_), .B2(G197gat), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n369_), .A2(KEYINPUT86), .A3(new_n370_), .A4(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n359_), .A3(G204gat), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n371_), .A2(new_n374_), .A3(new_n370_), .A4(new_n362_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n366_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n371_), .A2(new_n374_), .A3(new_n362_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n365_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT21), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n358_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G78gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n366_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n375_), .A2(new_n376_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n375_), .A2(new_n376_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n381_), .ZN(new_n389_));
  INV_X1    g188(.A(G78gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n358_), .ZN(new_n391_));
  AND2_X1   g190(.A1(G228gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT87), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n389_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n262_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n395_), .A2(new_n262_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n384_), .B(new_n391_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n398_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n384_), .A2(new_n391_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n396_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G22gat), .B(G50gat), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n353_), .A2(new_n357_), .A3(KEYINPUT29), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT28), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n406_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n404_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n409_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n404_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n411_), .A2(new_n407_), .A3(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT88), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n410_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n413_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n403_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n403_), .A2(new_n414_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G183gat), .A2(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT23), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT23), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(G183gat), .A3(G190gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G183gat), .ZN(new_n428_));
  INV_X1    g227(.A(G190gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT90), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT22), .ZN(new_n436_));
  INV_X1    g235(.A(G169gat), .ZN(new_n437_));
  INV_X1    g236(.A(G176gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n432_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n431_), .A2(new_n435_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT24), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(G169gat), .B2(G176gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G169gat), .A2(G176gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT80), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(G169gat), .B2(G176gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT25), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G183gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n428_), .A2(KEYINPUT25), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n429_), .A2(KEYINPUT26), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT26), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G190gat), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .A4(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n445_), .A2(new_n443_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n449_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n424_), .A2(new_n426_), .A3(KEYINPUT82), .ZN(new_n459_));
  OR3_X1    g258(.A1(new_n423_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n442_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT91), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n446_), .A2(new_n448_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n466_), .B(new_n427_), .C1(new_n467_), .C2(KEYINPUT24), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT24), .B1(new_n446_), .B2(new_n448_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n427_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT81), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n453_), .A2(new_n455_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT79), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n451_), .A2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n451_), .A2(new_n452_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n472_), .B(new_n474_), .C1(new_n475_), .C2(new_n473_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n468_), .A2(new_n471_), .A3(new_n476_), .A4(new_n449_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n459_), .A2(new_n460_), .A3(new_n430_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n459_), .A2(new_n460_), .A3(KEYINPUT83), .A4(new_n430_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n433_), .A2(new_n434_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n477_), .A2(new_n483_), .A3(new_n388_), .A4(new_n381_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n462_), .B(KEYINPUT91), .C1(new_n378_), .C2(new_n382_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n465_), .A2(KEYINPUT20), .A3(new_n484_), .A4(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G226gat), .A2(G233gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT19), .Z(new_n488_));
  XOR2_X1   g287(.A(new_n488_), .B(KEYINPUT89), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT20), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n378_), .A2(new_n382_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n462_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n477_), .A2(new_n483_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n389_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n496_), .A3(new_n488_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G8gat), .B(G36gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT18), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G64gat), .B(G92gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  NAND3_X1  g300(.A1(new_n490_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT92), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n490_), .A2(new_n504_), .A3(new_n497_), .A4(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n490_), .A2(new_n497_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n501_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT27), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n494_), .A2(new_n496_), .ZN(new_n512_));
  OAI22_X1  g311(.A1(new_n512_), .A2(new_n488_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n507_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT27), .A3(new_n502_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n422_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G127gat), .B(G134gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G113gat), .B(G120gat), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n518_), .A2(new_n519_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n523_));
  NOR4_X1   g322(.A1(new_n341_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT84), .B1(new_n343_), .B2(new_n337_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n335_), .B1(new_n526_), .B2(new_n351_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n355_), .A2(new_n356_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n354_), .A2(new_n343_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n518_), .B(new_n519_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n523_), .A2(new_n532_), .A3(KEYINPUT4), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G225gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n523_), .B2(KEYINPUT4), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT93), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n523_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n523_), .A2(new_n532_), .A3(KEYINPUT96), .A4(new_n534_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n531_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n534_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n523_), .A2(new_n532_), .A3(KEYINPUT4), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n537_), .A2(new_n542_), .A3(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT95), .ZN(new_n551_));
  XOR2_X1   g350(.A(G1gat), .B(G29gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G57gat), .B(G85gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n551_), .A2(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n552_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n554_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n549_), .A2(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n537_), .A2(new_n542_), .A3(new_n560_), .A4(new_n548_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G71gat), .B(G99gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G43gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n495_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(new_n522_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G227gat), .A2(G233gat), .ZN(new_n570_));
  INV_X1    g369(.A(G15gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT30), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT31), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n569_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n517_), .A2(new_n565_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT97), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n534_), .B1(new_n523_), .B2(KEYINPUT4), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n533_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n523_), .A2(new_n532_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n534_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n560_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n563_), .A2(KEYINPUT33), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n563_), .A2(KEYINPUT33), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n578_), .B1(new_n587_), .B2(new_n509_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n537_), .A2(new_n548_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n560_), .A4(new_n542_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n563_), .A2(KEYINPUT33), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n583_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n501_), .B1(new_n490_), .B2(new_n497_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(KEYINPUT92), .B2(new_n502_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n593_), .A2(new_n595_), .A3(KEYINPUT97), .A4(new_n505_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n501_), .A2(KEYINPUT32), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n490_), .A2(new_n497_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT98), .ZN(new_n599_));
  INV_X1    g398(.A(new_n597_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n513_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n513_), .B2(new_n600_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n564_), .B(new_n598_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n588_), .A2(new_n596_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n422_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n516_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n420_), .A2(new_n421_), .A3(new_n564_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n604_), .A2(new_n605_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n577_), .B1(new_n608_), .B2(new_n576_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n236_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n311_), .A2(new_n246_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT34), .Z(new_n618_));
  INV_X1    g417(.A(KEYINPUT35), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT75), .Z(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n619_), .B2(new_n618_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n615_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT76), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT76), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n615_), .A2(new_n616_), .A3(new_n625_), .A4(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n310_), .A2(new_n274_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n620_), .B1(new_n628_), .B2(new_n614_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT72), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT72), .B(new_n620_), .C1(new_n628_), .C2(new_n614_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n613_), .B1(new_n627_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n627_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n627_), .A2(new_n633_), .A3(new_n637_), .A4(new_n635_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n634_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n609_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n331_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n202_), .B1(new_n644_), .B2(new_n564_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n609_), .A2(new_n256_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT37), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n641_), .A2(new_n647_), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT37), .B(new_n634_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AND4_X1   g449(.A1(new_n329_), .A2(new_n646_), .A3(new_n229_), .A4(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n564_), .B(KEYINPUT99), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n202_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT38), .B1(new_n645_), .B2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n655_), .B1(KEYINPUT38), .B2(new_n654_), .ZN(G1324gat));
  NAND3_X1  g455(.A1(new_n651_), .A2(new_n214_), .A3(new_n516_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n643_), .A2(new_n606_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(KEYINPUT101), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n214_), .B1(new_n658_), .B2(KEYINPUT101), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n659_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n657_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(G1325gat));
  OAI21_X1  g465(.A(G15gat), .B1(new_n643_), .B2(new_n575_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT41), .Z(new_n668_));
  NAND3_X1  g467(.A1(new_n651_), .A2(new_n571_), .A3(new_n576_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1326gat));
  XNOR2_X1  g469(.A(new_n422_), .B(KEYINPUT102), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G22gat), .B1(new_n643_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT42), .ZN(new_n674_));
  INV_X1    g473(.A(G22gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n651_), .A2(new_n675_), .A3(new_n671_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1327gat));
  INV_X1    g476(.A(new_n641_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n646_), .A2(new_n678_), .A3(new_n329_), .A4(new_n228_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT105), .Z(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n564_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n650_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n609_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n604_), .A2(new_n605_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n606_), .A2(new_n607_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n576_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NOR4_X1   g486(.A1(new_n422_), .A2(new_n516_), .A3(new_n564_), .A4(new_n575_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT103), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n690_), .B(new_n577_), .C1(new_n608_), .C2(new_n576_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n689_), .A2(new_n682_), .A3(new_n691_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n692_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT104), .B1(new_n692_), .B2(KEYINPUT43), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n684_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n256_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n329_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n229_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT44), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n652_), .A2(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n681_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n699_), .B(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G36gat), .B1(new_n704_), .B2(new_n606_), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n516_), .A2(KEYINPUT106), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n516_), .A2(KEYINPUT106), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n680_), .A2(new_n706_), .A3(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT45), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n705_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n705_), .A2(KEYINPUT46), .A3(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  NAND3_X1  g515(.A1(new_n700_), .A2(G43gat), .A3(new_n576_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n680_), .A2(new_n576_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n718_), .A2(G43gat), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT47), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n717_), .A2(new_n722_), .A3(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1330gat));
  OAI21_X1  g523(.A(G50gat), .B1(new_n704_), .B2(new_n605_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n672_), .A2(G50gat), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT107), .Z(new_n727_));
  NAND2_X1  g526(.A1(new_n680_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT108), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n725_), .A2(new_n731_), .A3(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1331gat));
  NOR3_X1   g532(.A1(new_n228_), .A2(new_n256_), .A3(new_n329_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n642_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n565_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n609_), .A2(new_n696_), .ZN(new_n738_));
  AND4_X1   g537(.A1(new_n697_), .A2(new_n738_), .A3(new_n229_), .A4(new_n650_), .ZN(new_n739_));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n652_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n735_), .B2(new_n709_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT48), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n739_), .A2(new_n743_), .A3(new_n709_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1333gat));
  INV_X1    g546(.A(G71gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n735_), .B2(new_n576_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n739_), .A2(new_n748_), .A3(new_n576_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT110), .Z(G1334gat));
  AOI21_X1  g553(.A(new_n390_), .B1(new_n735_), .B2(new_n671_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT50), .Z(new_n756_));
  NAND3_X1  g555(.A1(new_n739_), .A2(new_n390_), .A3(new_n671_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT111), .Z(G1335gat));
  NAND4_X1  g558(.A1(new_n738_), .A2(new_n678_), .A3(new_n697_), .A4(new_n228_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n265_), .A3(new_n652_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT112), .B(new_n684_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n228_), .A2(new_n697_), .A3(new_n696_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT113), .Z(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n692_), .A2(KEYINPUT43), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n692_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT112), .B1(new_n771_), .B2(new_n684_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT114), .B1(new_n766_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n695_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n765_), .A4(new_n763_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n773_), .A2(new_n564_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n762_), .B1(new_n778_), .B2(new_n265_), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n761_), .A2(new_n266_), .A3(new_n516_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n773_), .A2(new_n709_), .A3(new_n777_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n266_), .ZN(G1337gat));
  NAND3_X1  g581(.A1(new_n773_), .A2(new_n576_), .A3(new_n777_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G99gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n761_), .A2(new_n576_), .A3(new_n263_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT51), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(new_n788_), .A3(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1338gat));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  OAI21_X1  g590(.A(G106gat), .B1(new_n791_), .B2(KEYINPUT115), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n765_), .A2(new_n422_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n695_), .B2(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n791_), .A2(KEYINPUT115), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n761_), .A2(new_n262_), .A3(new_n422_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n228_), .A2(new_n256_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n329_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT116), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n803_), .A3(new_n329_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n682_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT54), .ZN(new_n806_));
  INV_X1    g605(.A(new_n251_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n247_), .A2(new_n249_), .A3(new_n239_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n254_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n807_), .A2(new_n254_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n696_), .A2(new_n322_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n315_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT117), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n315_), .A2(new_n816_), .A3(new_n813_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n295_), .A2(new_n209_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n818_), .A2(KEYINPUT55), .A3(new_n300_), .A4(new_n304_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n304_), .A2(new_n314_), .A3(new_n296_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n301_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n815_), .A2(new_n817_), .A3(new_n819_), .A4(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT118), .B1(new_n822_), .B2(new_n319_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n812_), .B1(new_n823_), .B2(KEYINPUT56), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n821_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n816_), .B1(new_n315_), .B2(new_n813_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n320_), .B1(new_n827_), .B2(new_n817_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n828_), .A2(KEYINPUT118), .A3(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n811_), .B1(new_n824_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n641_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT119), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n828_), .B2(KEYINPUT118), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n822_), .A2(new_n319_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(KEYINPUT56), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n837_), .A3(new_n812_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n678_), .B1(new_n838_), .B2(new_n811_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n833_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n832_), .A2(new_n842_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n828_), .A2(new_n829_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n835_), .A2(KEYINPUT56), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n810_), .A2(new_n321_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n850_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n682_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n843_), .A2(new_n845_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n229_), .B1(new_n854_), .B2(KEYINPUT121), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n843_), .A2(new_n845_), .A3(new_n856_), .A4(new_n853_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n806_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n517_), .A2(new_n576_), .A3(new_n652_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT59), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n842_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n861_));
  AOI211_X1 g660(.A(KEYINPUT119), .B(new_n678_), .C1(new_n838_), .C2(new_n811_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n853_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n843_), .A2(KEYINPUT122), .A3(new_n853_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n845_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n228_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n806_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n859_), .A2(KEYINPUT59), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n860_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G113gat), .B1(new_n873_), .B2(new_n696_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n854_), .A2(KEYINPUT121), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n228_), .A3(new_n857_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n869_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n859_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n696_), .A2(G113gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n874_), .B1(new_n879_), .B2(new_n880_), .ZN(G1340gat));
  OAI21_X1  g680(.A(G120gat), .B1(new_n873_), .B2(new_n329_), .ZN(new_n882_));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n329_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(KEYINPUT60), .B2(new_n883_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n882_), .B1(new_n879_), .B2(new_n885_), .ZN(G1341gat));
  OAI21_X1  g685(.A(G127gat), .B1(new_n873_), .B2(new_n228_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n228_), .A2(G127gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n879_), .B2(new_n888_), .ZN(G1342gat));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n650_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n860_), .A2(new_n872_), .A3(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n879_), .B2(new_n641_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT123), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n892_), .A2(new_n893_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1343gat));
  INV_X1    g697(.A(new_n709_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n605_), .A2(new_n576_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n877_), .A2(new_n652_), .A3(new_n899_), .A4(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n696_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT124), .B(G141gat), .Z(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1344gat));
  NOR2_X1   g703(.A1(new_n901_), .A2(new_n329_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n339_), .ZN(G1345gat));
  NOR2_X1   g705(.A1(new_n901_), .A2(new_n228_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT61), .B(G155gat), .Z(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n901_), .B2(new_n650_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n641_), .A2(G162gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n901_), .B2(new_n911_), .ZN(G1347gat));
  NOR3_X1   g711(.A1(new_n899_), .A2(new_n575_), .A3(new_n652_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n870_), .A2(new_n256_), .A3(new_n672_), .A4(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT62), .B(new_n437_), .C1(new_n914_), .C2(KEYINPUT22), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n806_), .B1(new_n867_), .B2(new_n228_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n913_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n917_), .A2(new_n696_), .A3(new_n671_), .A4(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n916_), .B1(new_n919_), .B2(new_n436_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G169gat), .B1(new_n914_), .B2(KEYINPUT62), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n915_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(G1348gat));
  NAND2_X1  g722(.A1(new_n877_), .A2(new_n605_), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n924_), .A2(new_n438_), .A3(new_n329_), .A4(new_n918_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n870_), .A2(new_n672_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n918_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n697_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n925_), .B1(new_n928_), .B2(new_n438_), .ZN(G1349gat));
  NAND2_X1  g728(.A1(new_n913_), .A2(new_n229_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n926_), .A2(new_n475_), .A3(new_n930_), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n924_), .A2(new_n930_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n428_), .B2(new_n932_), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n927_), .A2(new_n472_), .A3(new_n678_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n926_), .A2(new_n650_), .A3(new_n918_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n429_), .ZN(G1351gat));
  NAND2_X1  g735(.A1(new_n607_), .A2(new_n575_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT125), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n899_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n877_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n696_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT126), .B(G197gat), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n941_), .B(new_n942_), .ZN(G1352gat));
  NOR2_X1   g742(.A1(new_n940_), .A2(new_n329_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(new_n361_), .ZN(G1353gat));
  NOR2_X1   g744(.A1(new_n940_), .A2(new_n228_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  AND2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n946_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n949_), .B1(new_n946_), .B2(new_n947_), .ZN(G1354gat));
  XNOR2_X1  g749(.A(KEYINPUT127), .B(G218gat), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n940_), .A2(new_n650_), .A3(new_n951_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n877_), .A2(new_n678_), .A3(new_n939_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n952_), .B1(new_n953_), .B2(new_n951_), .ZN(G1355gat));
endmodule


