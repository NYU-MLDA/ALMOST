//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n208_), .B(new_n211_), .Z(new_n212_));
  NAND2_X1  g011(.A1(G229gat), .A2(G233gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT75), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n211_), .B(KEYINPUT15), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n208_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n208_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n211_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n221_), .A3(new_n213_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G113gat), .B(G141gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G169gat), .B(G197gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n224_), .B(new_n225_), .Z(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n217_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT76), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT83), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G141gat), .A2(G148gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT2), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n239_));
  OR2_X1    g038(.A1(G141gat), .A2(G148gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n238_), .B(new_n239_), .C1(new_n240_), .C2(KEYINPUT3), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n232_), .B(new_n233_), .C1(new_n235_), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(new_n232_), .B2(KEYINPUT1), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n232_), .A2(KEYINPUT1), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n233_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n232_), .A2(new_n244_), .A3(KEYINPUT1), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n240_), .B(new_n236_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n242_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT28), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(KEYINPUT28), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G22gat), .B(G50gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G78gat), .B(G106gat), .ZN(new_n259_));
  INV_X1    g058(.A(G233gat), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n260_), .A2(KEYINPUT84), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(KEYINPUT84), .ZN(new_n262_));
  OAI21_X1  g061(.A(G228gat), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT86), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT85), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT21), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n268_), .A2(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n272_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n266_), .A2(new_n274_), .A3(new_n270_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n242_), .A2(new_n249_), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n263_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n275_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n274_), .B1(new_n266_), .B2(new_n270_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n263_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n243_), .B1(new_n242_), .B2(new_n249_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT87), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n263_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT87), .ZN(new_n288_));
  INV_X1    g087(.A(new_n284_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  AOI211_X1 g089(.A(new_n259_), .B(new_n280_), .C1(new_n285_), .C2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n280_), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n283_), .A2(KEYINPUT87), .A3(new_n284_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n288_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n259_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT89), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n291_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n280_), .B1(new_n285_), .B2(new_n290_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n259_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n297_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n258_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT90), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n258_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n297_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n299_), .A2(new_n300_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n306_), .B1(new_n309_), .B2(new_n301_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT90), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n296_), .A2(KEYINPUT91), .ZN(new_n312_));
  OR3_X1    g111(.A1(new_n299_), .A2(KEYINPUT91), .A3(new_n300_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n291_), .A2(new_n258_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n305_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT19), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT23), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT25), .B(G183gat), .Z(new_n325_));
  INV_X1    g124(.A(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT26), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT26), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(G176gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n334_), .A2(new_n322_), .A3(new_n321_), .ZN(new_n335_));
  OR3_X1    g134(.A1(new_n324_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n320_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT22), .ZN(new_n339_));
  OR2_X1    g138(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT78), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(G169gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n333_), .B(new_n345_), .C1(new_n342_), .C2(KEYINPUT78), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n338_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n273_), .A2(new_n275_), .A3(new_n336_), .A4(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(KEYINPUT92), .A3(KEYINPUT20), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT94), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n334_), .B(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(new_n337_), .B2(new_n320_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n332_), .A2(KEYINPUT22), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n345_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT95), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n333_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n330_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n325_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n324_), .A2(new_n335_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n276_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n349_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT92), .B1(new_n348_), .B2(KEYINPUT20), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n318_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n357_), .A2(new_n363_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n281_), .A2(new_n282_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n318_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n336_), .A2(new_n347_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT96), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n276_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n375_), .B1(new_n276_), .B2(new_n374_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n372_), .B(new_n373_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n368_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT18), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n368_), .A2(new_n384_), .A3(new_n379_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n387_), .A2(KEYINPUT27), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n372_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT99), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n318_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT20), .B1(new_n364_), .B2(new_n276_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n276_), .A2(new_n374_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT96), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n395_), .B1(new_n397_), .B2(new_n376_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT99), .B1(new_n398_), .B2(new_n373_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n366_), .A2(new_n318_), .A3(new_n367_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n385_), .B(new_n394_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n391_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n390_), .A2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT100), .B1(new_n316_), .B2(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G127gat), .B(G134gat), .Z(new_n405_));
  XOR2_X1   g204(.A(G113gat), .B(G120gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n277_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n242_), .A3(new_n249_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n409_), .A2(KEYINPUT4), .A3(new_n410_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n277_), .A2(new_n408_), .A3(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n413_), .B1(new_n417_), .B2(new_n412_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G57gat), .B(G85gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n418_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426_));
  INV_X1    g225(.A(G43gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT79), .B(G15gat), .Z(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n374_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n435_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n432_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n436_), .B2(new_n432_), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n407_), .B(KEYINPUT31), .Z(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n441_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n313_), .A2(new_n314_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n303_), .A2(new_n304_), .B1(new_n445_), .B2(new_n312_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n389_), .A2(new_n388_), .B1(new_n391_), .B2(new_n401_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT100), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .A4(new_n311_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n404_), .A2(new_n425_), .A3(new_n444_), .A4(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n315_), .B1(new_n310_), .B2(KEYINPUT90), .ZN(new_n451_));
  AOI211_X1 g250(.A(new_n304_), .B(new_n306_), .C1(new_n309_), .C2(new_n301_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n447_), .B(new_n425_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n418_), .A2(KEYINPUT98), .A3(KEYINPUT33), .A4(new_n423_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT98), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n412_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n411_), .A2(new_n412_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n423_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n455_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n417_), .A2(new_n412_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n411_), .A2(new_n412_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(new_n423_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n458_), .A2(new_n459_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n461_), .A2(new_n387_), .A3(new_n386_), .A4(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n384_), .A2(KEYINPUT32), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n394_), .B(new_n468_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n368_), .A2(new_n379_), .A3(new_n467_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n424_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n446_), .A2(new_n472_), .A3(new_n311_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n453_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT81), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n444_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n442_), .A2(KEYINPUT81), .A3(new_n443_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n231_), .B1(new_n450_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G230gat), .A2(G233gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(G85gat), .B(G92gat), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT9), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT10), .B(G99gat), .ZN(new_n485_));
  OAI221_X1 g284(.A(new_n483_), .B1(KEYINPUT9), .B2(new_n484_), .C1(G106gat), .C2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT6), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT64), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n486_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n482_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n497_), .B1(new_n492_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n491_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT66), .B1(new_n499_), .B2(new_n500_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n488_), .A2(new_n490_), .A3(KEYINPUT65), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  INV_X1    g307(.A(G99gat), .ZN(new_n509_));
  INV_X1    g308(.A(G106gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT66), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n498_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .A4(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n495_), .B1(new_n514_), .B2(new_n482_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n503_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AOI211_X1 g316(.A(KEYINPUT67), .B(new_n495_), .C1(new_n514_), .C2(new_n482_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n494_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G71gat), .B(G78gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(G57gat), .B(G64gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(KEYINPUT11), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n521_), .A2(new_n523_), .A3(KEYINPUT11), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n521_), .B2(KEYINPUT11), .ZN(new_n525_));
  OR3_X1    g324(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n519_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n530_), .B(new_n494_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n481_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT64), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n491_), .B(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n496_), .B1(new_n534_), .B2(new_n501_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n514_), .A2(new_n482_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT8), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n537_), .B2(KEYINPUT67), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n515_), .A2(new_n516_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n493_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT12), .B1(new_n540_), .B2(new_n530_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n519_), .A2(new_n542_), .A3(new_n528_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n481_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n540_), .B2(new_n530_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n532_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G120gat), .B(G148gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT5), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G176gat), .B(G204gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT69), .B1(new_n547_), .B2(new_n552_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n482_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n511_), .A2(new_n512_), .A3(new_n498_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n512_), .B1(new_n511_), .B2(new_n498_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n488_), .A2(new_n490_), .A3(KEYINPUT65), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT65), .B1(new_n488_), .B2(new_n490_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n557_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT67), .B1(new_n564_), .B2(new_n495_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(new_n539_), .A3(new_n503_), .ZN(new_n566_));
  AOI211_X1 g365(.A(KEYINPUT12), .B(new_n530_), .C1(new_n566_), .C2(new_n494_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n542_), .B1(new_n519_), .B2(new_n528_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n546_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n532_), .ZN(new_n570_));
  AND4_X1   g369(.A1(KEYINPUT69), .A2(new_n569_), .A3(new_n570_), .A4(new_n552_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n554_), .B(new_n555_), .C1(new_n556_), .C2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n547_), .A2(new_n552_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n571_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n553_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT70), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(KEYINPUT13), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n572_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n208_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n528_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n583_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n583_), .A2(new_n589_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT73), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n540_), .A2(new_n211_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n519_), .A2(new_n218_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT71), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT71), .B1(new_n519_), .B2(new_n218_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n598_), .A2(new_n595_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT72), .ZN(new_n608_));
  XOR2_X1   g407(.A(G134gat), .B(G162gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n605_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n614_), .B(new_n599_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n606_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n610_), .B(KEYINPUT36), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n606_), .B2(new_n615_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT37), .B1(new_n616_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n606_), .A2(new_n615_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n617_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n606_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n580_), .A2(new_n594_), .A3(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT74), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT74), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n480_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n203_), .A3(new_n424_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT101), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n228_), .A2(new_n229_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n580_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n616_), .A2(new_n619_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n450_), .B2(new_n479_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n593_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n203_), .B1(new_n642_), .B2(new_n424_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n632_), .B2(new_n631_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n634_), .A2(new_n644_), .ZN(G1324gat));
  NAND3_X1  g444(.A1(new_n630_), .A2(new_n204_), .A3(new_n403_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G8gat), .B1(new_n641_), .B2(new_n447_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(KEYINPUT39), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(KEYINPUT39), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n646_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g450(.A(G15gat), .B1(new_n641_), .B2(new_n478_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT41), .Z(new_n653_));
  INV_X1    g452(.A(G15gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n478_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n630_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(G1326gat));
  INV_X1    g456(.A(G22gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n630_), .A2(new_n658_), .A3(new_n316_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n316_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G22gat), .B1(new_n641_), .B2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(KEYINPUT42), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(KEYINPUT42), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(G1327gat));
  INV_X1    g463(.A(new_n594_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n639_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n480_), .A2(new_n580_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(G29gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n424_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n450_), .A2(new_n479_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n626_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT43), .B(new_n626_), .C1(new_n450_), .C2(new_n479_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n677_), .A2(KEYINPUT44), .A3(new_n665_), .A4(new_n638_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n675_), .A2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n638_), .A2(new_n665_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n424_), .A3(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT103), .ZN(new_n684_));
  OAI21_X1  g483(.A(G29gat), .B1(new_n683_), .B2(KEYINPUT103), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n671_), .B1(new_n684_), .B2(new_n685_), .ZN(G1328gat));
  NOR2_X1   g485(.A1(new_n447_), .A2(G36gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n669_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT105), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n669_), .A2(new_n690_), .A3(new_n687_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n689_), .A2(KEYINPUT45), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT45), .B1(new_n689_), .B2(new_n691_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n678_), .A2(new_n682_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G36gat), .B1(new_n695_), .B2(new_n447_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n694_), .A2(new_n696_), .A3(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n444_), .A2(G43gat), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n669_), .A2(new_n655_), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n695_), .A2(new_n702_), .B1(G43gat), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g504(.A(G50gat), .B1(new_n695_), .B2(new_n660_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n660_), .A2(G50gat), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT106), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n669_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(G1331gat));
  NOR2_X1   g509(.A1(new_n580_), .A2(new_n635_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n673_), .A2(new_n711_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n712_), .A2(new_n665_), .A3(new_n674_), .ZN(new_n713_));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n424_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n580_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n640_), .A2(new_n231_), .A3(new_n594_), .A4(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n425_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n717_), .B2(new_n447_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n713_), .A2(new_n723_), .A3(new_n403_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1333gat));
  OAI21_X1  g524(.A(G71gat), .B1(new_n717_), .B2(new_n478_), .ZN(new_n726_));
  XOR2_X1   g525(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G71gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n713_), .A2(new_n729_), .A3(new_n655_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n717_), .B2(new_n660_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G78gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n713_), .A2(new_n735_), .A3(new_n316_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1335gat));
  NOR3_X1   g536(.A1(new_n580_), .A2(new_n635_), .A3(new_n594_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n677_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n425_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n712_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n668_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n425_), .A2(G85gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(G1336gat));
  OAI21_X1  g543(.A(G92gat), .B1(new_n739_), .B2(new_n447_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n447_), .A2(G92gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n742_), .B2(new_n746_), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n739_), .B2(new_n478_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n485_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n444_), .A2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n742_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g551(.A(new_n316_), .B(new_n738_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G106gat), .B1(new_n753_), .B2(new_n754_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT52), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n677_), .A2(KEYINPUT110), .A3(new_n316_), .A4(new_n738_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n753_), .A2(new_n754_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .A4(G106gat), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n757_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n741_), .A2(new_n510_), .A3(new_n316_), .A4(new_n668_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT53), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n766_), .A3(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1339gat));
  NAND4_X1  g567(.A1(new_n580_), .A2(new_n231_), .A3(new_n594_), .A4(new_n626_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n769_), .B(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n212_), .A2(new_n213_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n219_), .A2(new_n221_), .A3(new_n214_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n227_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n229_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n575_), .A2(new_n576_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n554_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n546_), .B(KEYINPUT55), .C1(new_n567_), .C2(new_n568_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n544_), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n546_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n569_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n531_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n545_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n781_), .A2(new_n782_), .A3(new_n784_), .A4(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n551_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n551_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(KEYINPUT113), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n551_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT113), .A3(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n635_), .B1(new_n556_), .B2(new_n571_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n778_), .B1(new_n790_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n639_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(KEYINPUT57), .A3(new_n798_), .ZN(new_n799_));
  XOR2_X1   g598(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n800_));
  NAND2_X1  g599(.A1(new_n791_), .A2(new_n792_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n551_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n794_), .B1(new_n789_), .B2(KEYINPUT113), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n777_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n800_), .B1(new_n806_), .B2(new_n639_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n775_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n626_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT58), .B(new_n808_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n799_), .A2(new_n807_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n593_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n771_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n404_), .A2(new_n424_), .A3(new_n444_), .A4(new_n449_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(G113gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n635_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT59), .B1(new_n816_), .B2(new_n817_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n817_), .A2(KEYINPUT59), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n804_), .A2(new_n805_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n639_), .B1(new_n824_), .B2(new_n778_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n825_), .A2(KEYINPUT57), .B1(new_n812_), .B2(new_n811_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n594_), .B1(new_n826_), .B2(new_n807_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n827_), .B2(new_n771_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n821_), .A2(new_n822_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n822_), .B1(new_n821_), .B2(new_n828_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n231_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n820_), .B1(new_n831_), .B2(new_n819_), .ZN(G1340gat));
  NAND3_X1  g631(.A1(new_n821_), .A2(new_n716_), .A3(new_n828_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G120gat), .ZN(new_n834_));
  INV_X1    g633(.A(new_n818_), .ZN(new_n835_));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n580_), .B2(KEYINPUT60), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(KEYINPUT60), .B2(new_n836_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n834_), .B1(new_n835_), .B2(new_n838_), .ZN(G1341gat));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT116), .B(G127gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n815_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n829_), .A2(new_n830_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G127gat), .B1(new_n818_), .B2(new_n594_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n840_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n830_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n821_), .A2(new_n822_), .A3(new_n828_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n842_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n845_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(KEYINPUT117), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n846_), .A2(new_n851_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n818_), .A2(new_n853_), .A3(new_n639_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n829_), .A2(new_n830_), .A3(new_n626_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n853_), .ZN(G1343gat));
  NAND4_X1  g655(.A1(new_n478_), .A2(new_n424_), .A3(new_n316_), .A4(new_n447_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n816_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n635_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n716_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n594_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  AOI21_X1  g664(.A(G162gat), .B1(new_n858_), .B2(new_n639_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n674_), .A2(G162gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT118), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n858_), .B2(new_n868_), .ZN(G1347gat));
  NAND2_X1  g668(.A1(new_n814_), .A2(new_n665_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n771_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n478_), .A2(new_n424_), .A3(new_n316_), .A4(new_n447_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G169gat), .B1(new_n874_), .B2(new_n230_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n872_), .A2(new_n355_), .A3(new_n635_), .A4(new_n873_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(KEYINPUT62), .A3(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n879_), .B(G169gat), .C1(new_n874_), .C2(new_n230_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n877_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n878_), .B1(new_n877_), .B2(new_n880_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1348gat));
  INV_X1    g682(.A(new_n816_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n884_), .A2(new_n873_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(G176gat), .A3(new_n716_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n886_), .A2(KEYINPUT120), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n333_), .B1(new_n874_), .B2(new_n580_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(KEYINPUT120), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(G1349gat));
  AOI21_X1  g689(.A(G183gat), .B1(new_n885_), .B2(new_n594_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n874_), .A2(new_n360_), .A3(new_n815_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n874_), .B2(new_n626_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n895_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n639_), .A2(new_n359_), .ZN(new_n898_));
  XOR2_X1   g697(.A(new_n898_), .B(KEYINPUT122), .Z(new_n899_));
  OAI22_X1  g698(.A1(new_n896_), .A2(new_n897_), .B1(new_n874_), .B2(new_n899_), .ZN(G1351gat));
  NOR2_X1   g699(.A1(new_n447_), .A2(new_n424_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n478_), .A2(new_n316_), .A3(new_n901_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n816_), .A2(new_n230_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(G197gat), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n904_), .A2(KEYINPUT123), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(KEYINPUT123), .ZN(new_n906_));
  OR3_X1    g705(.A1(new_n903_), .A2(KEYINPUT124), .A3(G197gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT124), .B1(new_n903_), .B2(G197gat), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n905_), .A2(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1352gat));
  NOR2_X1   g708(.A1(new_n816_), .A2(new_n902_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n580_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT126), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n912_), .B(new_n914_), .ZN(G1353gat));
  NAND2_X1  g714(.A1(new_n910_), .A2(new_n593_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  AND2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(new_n916_), .B2(new_n917_), .ZN(G1354gat));
  NAND2_X1  g719(.A1(new_n910_), .A2(new_n639_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT127), .B(G218gat), .Z(new_n922_));
  NOR2_X1   g721(.A1(new_n626_), .A2(new_n922_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n921_), .A2(new_n922_), .B1(new_n910_), .B2(new_n923_), .ZN(G1355gat));
endmodule


