//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G85gat), .B(G92gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .A4(new_n211_), .ZN(new_n212_));
  NOR3_X1   g011(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT64), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(KEYINPUT64), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n214_), .A2(new_n208_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n205_), .A2(new_n219_), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n217_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n218_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n212_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G29gat), .B(G36gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT15), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n226_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n228_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G232gat), .A2(G233gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT34), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT35), .Z(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT70), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(KEYINPUT35), .A3(new_n233_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(KEYINPUT70), .A3(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT36), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G190gat), .B(G218gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT69), .ZN(new_n242_));
  XOR2_X1   g041(.A(G134gat), .B(G162gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n239_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(KEYINPUT36), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n237_), .A2(new_n238_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n247_), .A2(KEYINPUT71), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(KEYINPUT71), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n245_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n251_), .B1(KEYINPUT37), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G127gat), .B(G155gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT16), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G183gat), .B(G211gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT17), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G57gat), .B(G64gat), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT11), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(KEYINPUT11), .ZN(new_n264_));
  XOR2_X1   g063(.A(G71gat), .B(G78gat), .Z(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n264_), .A2(new_n265_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT73), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G15gat), .B(G22gat), .ZN(new_n272_));
  INV_X1    g071(.A(G1gat), .ZN(new_n273_));
  INV_X1    g072(.A(G8gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT14), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G1gat), .B(G8gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n271_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n261_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n280_), .B2(new_n279_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT74), .B(KEYINPUT17), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n260_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT75), .Z(new_n285_));
  OR2_X1    g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n256_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT77), .ZN(new_n290_));
  INV_X1    g089(.A(new_n268_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n223_), .A2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n268_), .B(new_n212_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(G230gat), .A3(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G230gat), .A2(G233gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n292_), .A2(KEYINPUT12), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT12), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n223_), .B2(new_n291_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n298_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n296_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n295_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G120gat), .B(G148gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT5), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G176gat), .B(G204gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n310_));
  INV_X1    g109(.A(new_n308_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n295_), .B(new_n311_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n304_), .A2(KEYINPUT67), .A3(new_n308_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n313_), .A2(new_n314_), .B1(new_n315_), .B2(KEYINPUT13), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n316_), .A2(new_n315_), .A3(KEYINPUT13), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n315_), .B2(KEYINPUT13), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n290_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT87), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT87), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G155gat), .A3(G162gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT1), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(KEYINPUT88), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT88), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n332_), .B2(new_n327_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n325_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n331_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n329_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT89), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n336_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n337_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT90), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n338_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n338_), .B2(new_n346_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n340_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT91), .B1(new_n349_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n338_), .A2(new_n346_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT90), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n338_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(new_n353_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT91), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n355_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n325_), .A2(new_n328_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n344_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  AOI211_X1 g167(.A(KEYINPUT92), .B(new_n366_), .C1(new_n355_), .C2(new_n364_), .ZN(new_n369_));
  OAI22_X1  g168(.A1(new_n342_), .A2(new_n343_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT93), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n336_), .A2(new_n341_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT89), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n336_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT93), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n349_), .A2(new_n354_), .A3(KEYINPUT91), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n363_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n367_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT92), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n365_), .A2(new_n344_), .A3(new_n367_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n375_), .A2(new_n376_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n371_), .A2(KEYINPUT29), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G211gat), .B(G218gat), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT21), .ZN(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT95), .B(G197gat), .Z(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G204gat), .ZN(new_n388_));
  INV_X1    g187(.A(G204gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n391_));
  INV_X1    g190(.A(G197gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(G204gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n386_), .B1(new_n395_), .B2(KEYINPUT97), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT97), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT21), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n387_), .A2(new_n389_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(G197gat), .B2(G204gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n385_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n396_), .A2(new_n398_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(G228gat), .B2(G233gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n384_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(new_n375_), .B2(new_n382_), .ZN(new_n408_));
  OAI211_X1 g207(.A(G228gat), .B(G233gat), .C1(new_n408_), .C2(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n411_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n406_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT28), .B(G22gat), .ZN(new_n416_));
  INV_X1    g215(.A(G50gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT94), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n371_), .A2(new_n383_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(new_n407_), .ZN(new_n422_));
  AOI211_X1 g221(.A(KEYINPUT94), .B(KEYINPUT29), .C1(new_n371_), .C2(new_n383_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n370_), .A2(KEYINPUT93), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n376_), .B1(new_n375_), .B2(new_n382_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n407_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT94), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n421_), .A2(new_n420_), .A3(new_n407_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n418_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n415_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n412_), .A2(new_n424_), .A3(new_n430_), .A4(new_n414_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G127gat), .B(G134gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT85), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G113gat), .B(G120gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n439_), .B(KEYINPUT31), .Z(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(KEYINPUT84), .B(G43gat), .Z(new_n442_));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(KEYINPUT23), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(KEYINPUT23), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT23), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G183gat), .A3(G190gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n445_), .B1(new_n449_), .B2(new_n443_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT82), .B(G169gat), .ZN(new_n453_));
  INV_X1    g252(.A(G176gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT22), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n454_), .B1(new_n455_), .B2(KEYINPUT81), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n453_), .B(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G169gat), .A2(G176gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT24), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G169gat), .A2(G176gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT24), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G190gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT79), .A3(KEYINPUT26), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT79), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT26), .B(G190gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(G183gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT78), .B1(new_n474_), .B2(KEYINPUT25), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT25), .B(G183gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT78), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n467_), .B1(new_n473_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n449_), .B(new_n462_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT26), .B(G190gat), .Z(new_n483_));
  OAI21_X1  g282(.A(new_n469_), .B1(new_n483_), .B2(KEYINPUT79), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT25), .B(G183gat), .Z(new_n485_));
  AOI21_X1  g284(.A(new_n475_), .B1(new_n485_), .B2(KEYINPUT78), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT80), .B1(new_n487_), .B2(new_n467_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n459_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT30), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G99gat), .ZN(new_n492_));
  OAI211_X1 g291(.A(KEYINPUT30), .B(new_n459_), .C1(new_n482_), .C2(new_n488_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n442_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n449_), .A2(new_n462_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n484_), .A2(new_n486_), .B1(new_n466_), .B2(new_n465_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(KEYINPUT80), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n480_), .A2(new_n481_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n458_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(KEYINPUT30), .ZN(new_n502_));
  INV_X1    g301(.A(new_n493_), .ZN(new_n503_));
  OAI21_X1  g302(.A(G99gat), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n442_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(G15gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G71gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n496_), .A2(new_n507_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT86), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n496_), .B2(new_n507_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n441_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n496_), .A2(new_n507_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n511_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n518_), .A2(KEYINPUT86), .A3(new_n512_), .A4(new_n440_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT27), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n403_), .B1(new_n394_), .B2(KEYINPUT21), .ZN(new_n523_));
  OAI211_X1 g322(.A(KEYINPUT21), .B(new_n385_), .C1(new_n394_), .C2(new_n397_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n394_), .A2(new_n397_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT22), .B(G169gat), .Z(new_n527_));
  OAI21_X1  g326(.A(new_n463_), .B1(new_n527_), .B2(G176gat), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n451_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n462_), .B1(new_n485_), .B2(new_n483_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(new_n450_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT98), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n460_), .B1(new_n464_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n533_), .B2(new_n464_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n530_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n522_), .B1(new_n526_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n526_), .B2(new_n489_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G226gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT19), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n522_), .B1(new_n404_), .B2(new_n536_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n543_), .B(new_n544_), .C1(new_n404_), .C2(new_n501_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G8gat), .B(G36gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT18), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G64gat), .B(G92gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  AND3_X1   g348(.A1(new_n542_), .A2(new_n545_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n521_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n538_), .B(new_n544_), .C1(new_n526_), .C2(new_n489_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT20), .B1(new_n526_), .B2(new_n537_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n526_), .B2(new_n489_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n555_), .B2(new_n544_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n549_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n542_), .A2(new_n545_), .A3(new_n549_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(KEYINPUT27), .A3(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n552_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n435_), .A2(new_n520_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT104), .ZN(new_n563_));
  AND4_X1   g362(.A1(new_n430_), .A2(new_n412_), .A3(new_n424_), .A4(new_n414_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n414_), .A2(new_n412_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n563_), .B(new_n561_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n515_), .A2(new_n519_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n563_), .B1(new_n434_), .B2(new_n561_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n562_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n371_), .A2(new_n383_), .A3(new_n439_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n370_), .A2(new_n439_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(KEYINPUT4), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT99), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n571_), .A2(KEYINPUT99), .A3(KEYINPUT4), .A4(new_n572_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT4), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n371_), .A2(new_n383_), .A3(new_n578_), .A4(new_n439_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G225gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT100), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G1gat), .B(G29gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G85gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT0), .B(G57gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  INV_X1    g387(.A(new_n581_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n571_), .A2(new_n572_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT101), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n584_), .A2(new_n588_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n588_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT101), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n590_), .B(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n582_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n593_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n597_), .A3(KEYINPUT103), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n599_), .B(new_n593_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n549_), .A2(KEYINPUT32), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n542_), .A2(new_n545_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT102), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n556_), .A2(new_n602_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n603_), .A2(KEYINPUT102), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n605_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n598_), .A2(new_n600_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n592_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n550_), .A2(new_n551_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n584_), .A2(KEYINPUT33), .A3(new_n588_), .A4(new_n591_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n577_), .A2(new_n589_), .A3(new_n579_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n571_), .A2(new_n572_), .A3(new_n581_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n593_), .A3(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .A4(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n609_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n435_), .A2(new_n567_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n570_), .A2(new_n601_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n278_), .B(new_n226_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n278_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n227_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n278_), .B2(new_n226_), .ZN(new_n626_));
  AOI22_X1  g425(.A1(new_n621_), .A2(new_n623_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(G113gat), .B(G141gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(G169gat), .B(G197gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n627_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n620_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n320_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n601_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n273_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n248_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n620_), .A2(new_n638_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n319_), .A2(new_n287_), .A3(new_n632_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(new_n636_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n637_), .B1(new_n273_), .B2(new_n642_), .ZN(new_n643_));
  MUX2_X1   g442(.A(new_n637_), .B(new_n643_), .S(KEYINPUT38), .Z(G1324gat));
  INV_X1    g443(.A(new_n561_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n635_), .A2(new_n274_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(new_n645_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(KEYINPUT39), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n274_), .B1(new_n648_), .B2(KEYINPUT39), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n649_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n646_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1325gat));
  NAND2_X1  g455(.A1(new_n641_), .A2(new_n567_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G15gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n635_), .A2(new_n509_), .A3(new_n567_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n641_), .B2(new_n435_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n635_), .A2(new_n664_), .A3(new_n435_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1327gat));
  INV_X1    g468(.A(new_n319_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n287_), .A3(new_n631_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n570_), .A2(new_n601_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n618_), .A2(new_n619_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n673_), .B1(new_n676_), .B2(new_n255_), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT43), .B(new_n256_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n672_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n620_), .B2(new_n256_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n434_), .A2(new_n561_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT104), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n567_), .A3(new_n566_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n636_), .B1(new_n686_), .B2(new_n562_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n619_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n609_), .B2(new_n617_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n673_), .B(new_n255_), .C1(new_n687_), .C2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n671_), .B1(new_n683_), .B2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT108), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n682_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(KEYINPUT44), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n693_), .A2(G29gat), .A3(new_n636_), .A4(new_n694_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n319_), .A2(new_n248_), .A3(new_n288_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n633_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n636_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n695_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n695_), .A2(KEYINPUT109), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1328gat));
  XNOR2_X1  g504(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n561_), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n693_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n645_), .A2(new_n708_), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n697_), .A2(KEYINPUT45), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT45), .B1(new_n697_), .B2(new_n711_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n707_), .B1(new_n710_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n694_), .A2(new_n645_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n692_), .B2(new_n682_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n714_), .B(new_n706_), .C1(new_n718_), .C2(new_n708_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1329gat));
  NAND4_X1  g519(.A1(new_n693_), .A2(G43gat), .A3(new_n567_), .A4(new_n694_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G43gat), .B1(new_n698_), .B2(new_n567_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT47), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n721_), .A2(new_n726_), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1330gat));
  NAND3_X1  g527(.A1(new_n698_), .A2(new_n417_), .A3(new_n435_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n434_), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n693_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G50gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n693_), .B2(new_n730_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(G1331gat));
  NOR2_X1   g534(.A1(new_n287_), .A2(new_n631_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n639_), .A2(new_n319_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n601_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n676_), .A2(new_n632_), .ZN(new_n741_));
  OR4_X1    g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n290_), .A4(new_n670_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n290_), .A2(new_n670_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n743_), .B2(new_n741_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n738_), .B1(new_n745_), .B2(new_n601_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT113), .B(new_n738_), .C1(new_n745_), .C2(new_n601_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n739_), .B1(new_n748_), .B2(new_n749_), .ZN(G1332gat));
  OAI21_X1  g549(.A(G64gat), .B1(new_n737_), .B2(new_n561_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT114), .Z(new_n752_));
  OR2_X1    g551(.A1(new_n752_), .A2(KEYINPUT48), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(KEYINPUT48), .ZN(new_n754_));
  OR3_X1    g553(.A1(new_n745_), .A2(G64gat), .A3(new_n561_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n737_), .B2(new_n520_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n520_), .A2(G71gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n745_), .B2(new_n760_), .ZN(G1334gat));
  OAI21_X1  g560(.A(G78gat), .B1(new_n737_), .B2(new_n434_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT50), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n434_), .A2(G78gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n745_), .B2(new_n764_), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n677_), .A2(new_n678_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n319_), .A2(new_n287_), .A3(new_n632_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769_), .B2(new_n601_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n620_), .A2(new_n631_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n670_), .A2(new_n248_), .A3(new_n288_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n209_), .A3(new_n636_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n775_), .ZN(G1336gat));
  OAI21_X1  g575(.A(G92gat), .B1(new_n769_), .B2(new_n561_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n210_), .A3(new_n645_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1337gat));
  AND3_X1   g578(.A1(new_n774_), .A2(new_n567_), .A3(new_n202_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n768_), .A2(new_n567_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(G99gat), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT51), .Z(G1338gat));
  NOR3_X1   g582(.A1(new_n773_), .A2(G106gat), .A3(new_n434_), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n434_), .B(new_n767_), .C1(new_n683_), .C2(new_n690_), .ZN(new_n785_));
  OR3_X1    g584(.A1(new_n785_), .A2(KEYINPUT52), .A3(new_n203_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT52), .B1(new_n785_), .B2(new_n203_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n784_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n788_), .B(new_n790_), .ZN(G1339gat));
  NOR2_X1   g590(.A1(new_n686_), .A2(new_n601_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n299_), .A2(new_n301_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n303_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n794_), .A2(KEYINPUT55), .A3(new_n795_), .A4(new_n298_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n293_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(G230gat), .A3(G233gat), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n796_), .A2(new_n798_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n308_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n308_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n630_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n625_), .B(new_n623_), .C1(new_n229_), .C2(new_n624_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n627_), .A2(new_n630_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n312_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n806_), .A2(KEYINPUT58), .A3(new_n810_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n255_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n804_), .A2(new_n817_), .A3(new_n805_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n801_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n308_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n312_), .A2(new_n631_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n313_), .A2(new_n314_), .A3(new_n809_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n816_), .B1(new_n824_), .B2(new_n248_), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT57), .B(new_n638_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n815_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n288_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT118), .B(new_n815_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n256_), .A2(new_n736_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT54), .B1(new_n832_), .B2(new_n319_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n670_), .A2(new_n256_), .A3(new_n834_), .A4(new_n736_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n793_), .B1(new_n831_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n631_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n829_), .A2(new_n830_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT59), .B1(new_n840_), .B2(new_n793_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n827_), .A2(new_n287_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n836_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n792_), .A2(KEYINPUT119), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n792_), .A2(KEYINPUT119), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .A4(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n841_), .A2(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n848_), .A2(new_n631_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n839_), .B1(new_n849_), .B2(new_n838_), .ZN(G1340gat));
  OAI211_X1 g649(.A(new_n319_), .B(new_n847_), .C1(new_n837_), .C2(new_n844_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n670_), .B2(G120gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n837_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n841_), .A2(KEYINPUT120), .A3(new_n319_), .A4(new_n847_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n853_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G120gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n837_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1341gat));
  INV_X1    g660(.A(G127gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n837_), .A2(new_n862_), .A3(new_n288_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n848_), .A2(new_n288_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n837_), .A2(new_n866_), .A3(new_n638_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n848_), .A2(new_n255_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n866_), .ZN(G1343gat));
  NAND2_X1  g668(.A1(new_n831_), .A2(new_n836_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n562_), .A2(new_n601_), .ZN(new_n871_));
  XOR2_X1   g670(.A(new_n871_), .B(KEYINPUT121), .Z(new_n872_));
  AND2_X1   g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n631_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n319_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n873_), .A2(new_n878_), .A3(new_n288_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n870_), .A2(new_n872_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT122), .B1(new_n880_), .B2(new_n287_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n882_), .B(new_n884_), .ZN(G1346gat));
  OR3_X1    g684(.A1(new_n880_), .A2(G162gat), .A3(new_n248_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G162gat), .B1(new_n880_), .B2(new_n256_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1347gat));
  AOI21_X1  g687(.A(new_n435_), .B1(new_n836_), .B2(new_n842_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n636_), .A2(new_n520_), .A3(new_n561_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n631_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G169gat), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(KEYINPUT123), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(KEYINPUT123), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n893_), .A2(KEYINPUT62), .A3(new_n894_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n891_), .A2(new_n527_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(G1348gat));
  NAND2_X1  g699(.A1(new_n889_), .A2(new_n890_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G176gat), .B1(new_n902_), .B2(new_n319_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n840_), .A2(new_n435_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n890_), .A2(G176gat), .A3(new_n319_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  AND2_X1   g705(.A1(new_n890_), .A2(new_n288_), .ZN(new_n907_));
  AOI21_X1  g706(.A(G183gat), .B1(new_n904_), .B2(new_n907_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n907_), .A2(new_n485_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n889_), .B2(new_n909_), .ZN(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n901_), .B2(new_n256_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n638_), .A2(new_n472_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n901_), .B2(new_n912_), .ZN(G1351gat));
  NOR4_X1   g712(.A1(new_n636_), .A2(new_n434_), .A3(new_n567_), .A4(new_n561_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n870_), .A2(new_n914_), .ZN(new_n915_));
  OR4_X1    g714(.A1(KEYINPUT124), .A2(new_n915_), .A3(new_n392_), .A4(new_n632_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n870_), .A2(new_n914_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n631_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT124), .B1(new_n918_), .B2(new_n392_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n392_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n916_), .A2(new_n919_), .A3(new_n920_), .ZN(G1352gat));
  AOI21_X1  g720(.A(new_n670_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n917_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n923_), .B(new_n924_), .Z(G1353gat));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n915_), .B2(new_n287_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n928_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n915_), .A2(new_n287_), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT63), .B(G211gat), .Z(new_n932_));
  AOI22_X1  g731(.A1(new_n929_), .A2(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1354gat));
  INV_X1    g732(.A(G218gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n917_), .A2(new_n934_), .A3(new_n638_), .ZN(new_n935_));
  OAI21_X1  g734(.A(G218gat), .B1(new_n915_), .B2(new_n256_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n937_), .B(new_n938_), .ZN(G1355gat));
endmodule


