//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT64), .Z(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT6), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT10), .B(G99gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G106gat), .ZN(new_n208_));
  OAI221_X1 g007(.A(new_n205_), .B1(KEYINPUT9), .B2(new_n206_), .C1(new_n207_), .C2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G85gat), .B(G92gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT9), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(KEYINPUT66), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214_));
  INV_X1    g013(.A(new_n212_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n214_), .B1(new_n209_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n205_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(KEYINPUT8), .B(new_n211_), .C1(new_n218_), .C2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n211_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n213_), .A2(new_n216_), .A3(new_n222_), .A4(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G57gat), .B(G64gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT11), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(KEYINPUT11), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G71gat), .B(G78gat), .ZN(new_n230_));
  MUX2_X1   g029(.A(new_n228_), .B(new_n229_), .S(new_n230_), .Z(new_n231_));
  OR2_X1    g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n226_), .A2(new_n231_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n203_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(KEYINPUT12), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n203_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT68), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n238_), .B(new_n203_), .C1(new_n226_), .C2(new_n231_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT69), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(new_n240_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n234_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G120gat), .B(G148gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G204gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT5), .B(G176gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n249_), .B(KEYINPUT70), .Z(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n245_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT13), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT13), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n251_), .B(new_n255_), .C1(new_n245_), .C2(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G43gat), .B(G50gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(G29gat), .B(G36gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT15), .Z(new_n263_));
  XNOR2_X1  g062(.A(G15gat), .B(G22gat), .ZN(new_n264_));
  INV_X1    g063(.A(G1gat), .ZN(new_n265_));
  INV_X1    g064(.A(G8gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT14), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G1gat), .B(G8gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n263_), .A2(KEYINPUT75), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(new_n262_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT75), .B1(new_n263_), .B2(new_n270_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G229gat), .A2(G233gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n270_), .B(new_n262_), .Z(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G113gat), .B(G141gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G169gat), .B(G197gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n279_), .B(new_n282_), .Z(new_n283_));
  NOR2_X1   g082(.A1(new_n259_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT107), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT20), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT91), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT90), .B(G204gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(G197gat), .ZN(new_n289_));
  INV_X1    g088(.A(G204gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G197gat), .ZN(new_n291_));
  OR2_X1    g090(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n292_));
  INV_X1    g091(.A(G197gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n292_), .A2(KEYINPUT91), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n291_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT21), .ZN(new_n297_));
  XOR2_X1   g096(.A(G211gat), .B(G218gat), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n293_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n290_), .A2(G197gat), .ZN(new_n301_));
  OR3_X1    g100(.A1(new_n300_), .A2(KEYINPUT21), .A3(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(KEYINPUT21), .B(new_n298_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT92), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT23), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G183gat), .A3(G190gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n315_), .A3(KEYINPUT79), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n317_), .A3(KEYINPUT23), .ZN(new_n318_));
  INV_X1    g117(.A(G183gat), .ZN(new_n319_));
  INV_X1    g118(.A(G190gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n316_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(G176gat), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT78), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n325_), .A2(KEYINPUT78), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n311_), .B(new_n322_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n313_), .A2(new_n315_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(KEYINPUT26), .B2(new_n320_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n320_), .A2(KEYINPUT26), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT26), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n337_), .B2(new_n332_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT25), .B(G183gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n331_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT24), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n310_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n340_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n329_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n286_), .B1(new_n307_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT19), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n325_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(KEYINPUT98), .A3(new_n311_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n330_), .A2(new_n321_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT98), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n325_), .B2(new_n310_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT99), .ZN(new_n362_));
  INV_X1    g161(.A(new_n337_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n339_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n349_), .A2(new_n364_), .A3(new_n318_), .A4(new_n316_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n357_), .A2(new_n360_), .A3(new_n366_), .A4(new_n358_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n352_), .B(new_n355_), .C1(new_n307_), .C2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n322_), .A2(new_n311_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n325_), .B(KEYINPUT78), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n370_), .A2(new_n371_), .B1(new_n340_), .B2(new_n349_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n373_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT97), .B1(new_n373_), .B2(KEYINPUT20), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n368_), .A2(new_n307_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n369_), .B1(new_n377_), .B2(new_n355_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G8gat), .B(G36gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n369_), .B(new_n385_), .C1(new_n377_), .C2(new_n355_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n373_), .A2(KEYINPUT20), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT97), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n368_), .A2(new_n307_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n373_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n392_), .A2(new_n355_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n303_), .A2(new_n306_), .A3(new_n365_), .A4(new_n361_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n352_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n354_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n383_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n386_), .A3(KEYINPUT27), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n389_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT1), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n405_));
  OR2_X1    g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n403_), .A2(KEYINPUT1), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT84), .B1(new_n410_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT1), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(G155gat), .B2(G162gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT83), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n409_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n404_), .A2(new_n406_), .A3(new_n405_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n423_));
  INV_X1    g222(.A(new_n414_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n415_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n406_), .A2(new_n403_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT86), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n406_), .A2(new_n429_), .A3(new_n403_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n413_), .A2(KEYINPUT2), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT2), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(G141gat), .A3(G148gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438_));
  INV_X1    g237(.A(G141gat), .ZN(new_n439_));
  INV_X1    g238(.A(G148gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(KEYINPUT85), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n441_), .A2(new_n437_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(new_n436_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n432_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT87), .B1(new_n426_), .B2(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n423_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n450_));
  OAI211_X1 g249(.A(KEYINPUT87), .B(new_n447_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT29), .B1(new_n448_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G228gat), .A2(G233gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT88), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT89), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n307_), .A3(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G78gat), .B(G106gat), .Z(new_n458_));
  NAND2_X1  g257(.A1(new_n442_), .A2(KEYINPUT85), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n445_), .A2(new_n444_), .A3(new_n436_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n431_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n415_), .B2(new_n425_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT93), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n447_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT29), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n307_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n455_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n457_), .A2(new_n458_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n458_), .B1(new_n457_), .B2(new_n469_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n465_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n463_), .A3(new_n451_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G50gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT28), .B(G22gat), .ZN(new_n476_));
  INV_X1    g275(.A(G50gat), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n473_), .A2(new_n463_), .A3(new_n477_), .A4(new_n451_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n475_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n476_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n480_));
  OAI22_X1  g279(.A1(new_n470_), .A2(new_n471_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT94), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n457_), .A2(new_n469_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n458_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n457_), .A2(new_n469_), .A3(new_n458_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n479_), .A2(new_n480_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT94), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n483_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n471_), .B(KEYINPUT95), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n479_), .A2(new_n480_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT96), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n487_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n457_), .A2(new_n469_), .A3(KEYINPUT96), .A4(new_n458_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n492_), .A2(new_n493_), .A3(new_n495_), .A4(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n402_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G113gat), .B(G120gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(G127gat), .B(G134gat), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n500_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G225gat), .A2(G233gat), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n503_), .A2(KEYINPUT101), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n503_), .A2(KEYINPUT101), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n465_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n503_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n473_), .B2(new_n451_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n508_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n513_), .B(new_n503_), .C1(new_n448_), .C2(new_n452_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n505_), .B(KEYINPUT102), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n510_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT103), .B(KEYINPUT0), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G85gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G1gat), .B(G29gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n510_), .B(new_n523_), .C1(new_n514_), .C2(new_n517_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n378_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n385_), .A2(KEYINPUT32), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT106), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n527_), .A2(new_n531_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n504_), .A2(new_n509_), .A3(new_n516_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n515_), .A2(new_n505_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n524_), .B(new_n537_), .C1(new_n514_), .C2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n384_), .A2(new_n386_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n526_), .A2(KEYINPUT105), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(KEYINPUT104), .A3(KEYINPUT33), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT104), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n526_), .B2(KEYINPUT105), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n526_), .B2(new_n544_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n536_), .B1(new_n543_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n481_), .A2(new_n482_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT94), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n493_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n471_), .B(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n550_), .B(new_n551_), .C1(new_n552_), .C2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n498_), .A2(new_n528_), .B1(new_n549_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n351_), .B(KEYINPUT30), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G227gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT80), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G71gat), .B(G99gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(KEYINPUT81), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G43gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n562_), .B1(new_n558_), .B2(KEYINPUT81), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n564_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n568_), .B(new_n569_), .C1(KEYINPUT81), .C2(new_n558_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT82), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n503_), .B(KEYINPUT31), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n572_), .B(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n285_), .B1(new_n557_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n402_), .A2(KEYINPUT108), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT27), .B1(new_n384_), .B2(new_n386_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n400_), .A2(new_n386_), .A3(KEYINPUT27), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT108), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n556_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n575_), .A2(new_n528_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n555_), .A2(new_n528_), .A3(new_n580_), .ZN(new_n587_));
  AOI211_X1 g386(.A(new_n544_), .B(new_n546_), .C1(new_n526_), .C2(KEYINPUT105), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n384_), .A2(new_n386_), .A3(new_n539_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n545_), .A2(new_n547_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n525_), .A2(new_n526_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n534_), .A2(new_n535_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n590_), .A2(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n587_), .B1(new_n594_), .B2(new_n555_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n575_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(KEYINPUT107), .A3(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n576_), .A2(new_n586_), .A3(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n284_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n226_), .A2(new_n262_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT73), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n604_));
  NAND2_X1  g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(KEYINPUT35), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n226_), .A2(new_n263_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n602_), .B(new_n608_), .C1(KEYINPUT35), .C2(new_n606_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n607_), .A2(new_n609_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT36), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n611_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n607_), .A2(new_n609_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(new_n610_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n601_), .B1(new_n617_), .B2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n619_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n616_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(new_n625_), .A3(new_n610_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n626_), .A3(new_n600_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n231_), .B(new_n270_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n628_), .B(new_n629_), .Z(new_n630_));
  INV_X1    g429(.A(KEYINPUT17), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G127gat), .B(G155gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(G211gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT16), .B(G183gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n630_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(KEYINPUT17), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n630_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n623_), .A2(new_n627_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n599_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT109), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n265_), .A3(new_n527_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT38), .ZN(new_n645_));
  INV_X1    g444(.A(new_n639_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n624_), .A2(new_n626_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n599_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n528_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(new_n650_), .ZN(G1324gat));
  OAI21_X1  g450(.A(G8gat), .B1(new_n649_), .B2(new_n583_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(new_n583_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n643_), .A2(new_n266_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n649_), .B2(new_n596_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT41), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n641_), .A2(G15gat), .A3(new_n596_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1326gat));
  OAI21_X1  g461(.A(G22gat), .B1(new_n649_), .B2(new_n556_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT42), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n556_), .A2(G22gat), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT110), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n599_), .A2(new_n640_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT111), .ZN(G1327gat));
  AND3_X1   g468(.A1(new_n595_), .A2(KEYINPUT107), .A3(new_n596_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT107), .B1(new_n595_), .B2(new_n596_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n584_), .A2(new_n585_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n647_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n284_), .A2(new_n646_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n527_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n623_), .A2(new_n627_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n598_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n598_), .B2(new_n681_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n646_), .B(new_n284_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n685_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n527_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n679_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  NAND3_X1  g489(.A1(new_n686_), .A2(new_n687_), .A3(new_n654_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n678_), .A2(new_n693_), .A3(new_n654_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT45), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n692_), .A2(new_n695_), .A3(KEYINPUT46), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  NAND3_X1  g499(.A1(new_n686_), .A2(new_n687_), .A3(new_n575_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n596_), .A2(G43gat), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n701_), .A2(G43gat), .B1(new_n678_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g503(.A1(new_n686_), .A2(new_n687_), .A3(new_n555_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT112), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(KEYINPUT112), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(G50gat), .A3(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n678_), .A2(new_n477_), .A3(new_n555_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1331gat));
  NAND2_X1  g509(.A1(new_n259_), .A2(new_n283_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n673_), .A2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n648_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(G57gat), .A3(new_n527_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n714_), .A2(KEYINPUT113), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(KEYINPUT113), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n712_), .A2(new_n640_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n528_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n715_), .B(new_n716_), .C1(G57gat), .C2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT114), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1332gat));
  INV_X1    g520(.A(G64gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n713_), .B2(new_n654_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT48), .Z(new_n724_));
  INV_X1    g523(.A(new_n717_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n722_), .A3(new_n654_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n713_), .B2(new_n575_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT49), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n728_), .A3(new_n575_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1334gat));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n713_), .B2(new_n555_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT50), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n725_), .A2(new_n733_), .A3(new_n555_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n711_), .A2(new_n639_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n675_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n527_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n681_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT43), .B1(new_n673_), .B2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n598_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n738_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n527_), .A2(G85gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n741_), .B1(new_n746_), .B2(new_n747_), .ZN(G1336gat));
  AOI21_X1  g547(.A(G92gat), .B1(new_n740_), .B2(new_n654_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n654_), .A2(G92gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n746_), .B2(new_n750_), .ZN(G1337gat));
  OR3_X1    g550(.A1(new_n739_), .A2(new_n207_), .A3(new_n596_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n746_), .A2(new_n575_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n753_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT115), .B1(new_n753_), .B2(G99gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT51), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n752_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1338gat));
  OAI211_X1 g559(.A(new_n555_), .B(new_n738_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT116), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n745_), .A2(new_n763_), .A3(new_n555_), .A4(new_n738_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n764_), .A3(G106gat), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT52), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n762_), .A2(new_n764_), .A3(new_n767_), .A4(G106gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  OR3_X1    g568(.A1(new_n739_), .A2(new_n208_), .A3(new_n556_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n769_), .A2(new_n773_), .A3(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  INV_X1    g574(.A(G113gat), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n235_), .A2(new_n232_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(new_n203_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n242_), .A2(new_n244_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n235_), .A2(new_n240_), .A3(KEYINPUT55), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n252_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT117), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n283_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n251_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n244_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n243_), .B1(new_n235_), .B2(new_n240_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n781_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n779_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n783_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n252_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n789_), .B1(new_n796_), .B2(new_n786_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n276_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n275_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n798_), .B2(new_n278_), .ZN(new_n800_));
  MUX2_X1   g599(.A(new_n279_), .B(new_n800_), .S(new_n282_), .Z(new_n801_));
  AOI22_X1  g600(.A1(new_n788_), .A2(new_n797_), .B1(new_n253_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n777_), .B1(new_n802_), .B2(new_n647_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n251_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n796_), .B2(KEYINPUT56), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n789_), .B1(new_n796_), .B2(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n784_), .A2(new_n785_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(KEYINPUT58), .A3(new_n809_), .A4(new_n801_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(new_n681_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n253_), .A2(new_n801_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n251_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n283_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n796_), .B2(new_n786_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n812_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(KEYINPUT57), .A3(new_n674_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n803_), .A2(new_n811_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n646_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n256_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n245_), .A2(new_n252_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n255_), .B1(new_n821_), .B2(new_n251_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n640_), .B(new_n283_), .C1(new_n820_), .C2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT118), .B1(new_n819_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n828_), .B(new_n825_), .C1(new_n818_), .C2(new_n646_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n584_), .A2(new_n596_), .A3(new_n528_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n776_), .B1(new_n832_), .B2(new_n283_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n833_), .A2(KEYINPUT119), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(KEYINPUT119), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n819_), .A2(new_n826_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(new_n831_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n832_), .B2(KEYINPUT59), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT121), .B(G113gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n814_), .A3(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n834_), .A2(new_n835_), .A3(new_n841_), .ZN(G1340gat));
  INV_X1    g641(.A(new_n832_), .ZN(new_n843_));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  INV_X1    g643(.A(new_n259_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(KEYINPUT60), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n844_), .A2(KEYINPUT60), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(KEYINPUT122), .B2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n843_), .B(new_n848_), .C1(KEYINPUT122), .C2(new_n846_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n839_), .A2(new_n259_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n844_), .ZN(G1341gat));
  AOI21_X1  g650(.A(G127gat), .B1(new_n843_), .B2(new_n639_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n639_), .A2(G127gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n839_), .B2(new_n853_), .ZN(G1342gat));
  AOI21_X1  g653(.A(G134gat), .B1(new_n843_), .B2(new_n647_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n681_), .A2(G134gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n839_), .B2(new_n856_), .ZN(G1343gat));
  NOR3_X1   g656(.A1(new_n827_), .A2(new_n829_), .A3(new_n575_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n858_), .A2(new_n527_), .A3(new_n583_), .A4(new_n555_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n283_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n439_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n845_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n440_), .ZN(G1345gat));
  NOR2_X1   g662(.A1(new_n859_), .A2(new_n646_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n864_), .B(new_n866_), .ZN(G1346gat));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n859_), .A2(new_n868_), .A3(new_n742_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n859_), .B2(new_n674_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT123), .B(new_n868_), .C1(new_n859_), .C2(new_n674_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n869_), .B1(new_n872_), .B2(new_n873_), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n583_), .A2(new_n527_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n575_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT124), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n814_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT125), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n555_), .B1(new_n819_), .B2(new_n826_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n308_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT62), .Z(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n877_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n323_), .A2(new_n324_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n814_), .A3(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n886_), .ZN(G1348gat));
  AOI21_X1  g686(.A(G176gat), .B1(new_n884_), .B2(new_n259_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n827_), .A2(new_n829_), .A3(new_n555_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n877_), .A2(G176gat), .A3(new_n259_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(G1349gat));
  NOR3_X1   g690(.A1(new_n883_), .A2(new_n646_), .A3(new_n339_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n639_), .A3(new_n877_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n319_), .ZN(G1350gat));
  OAI21_X1  g693(.A(G190gat), .B1(new_n883_), .B2(new_n742_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n647_), .A2(new_n363_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n883_), .B2(new_n896_), .ZN(G1351gat));
  NAND4_X1  g696(.A1(new_n830_), .A2(new_n555_), .A3(new_n596_), .A4(new_n875_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n283_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n293_), .ZN(G1352gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n845_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n288_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n290_), .B2(new_n901_), .ZN(G1353gat));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n904_));
  INV_X1    g703(.A(G211gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n836_), .A2(new_n828_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n819_), .A2(KEYINPUT118), .A3(new_n826_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n908_), .A2(new_n555_), .A3(new_n596_), .A4(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n875_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n910_), .A2(new_n646_), .A3(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n904_), .A2(new_n905_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n907_), .B1(new_n912_), .B2(new_n914_), .ZN(new_n915_));
  NOR4_X1   g714(.A1(new_n898_), .A2(KEYINPUT126), .A3(new_n646_), .A4(new_n913_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n906_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n912_), .A2(new_n907_), .A3(new_n914_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n858_), .A2(new_n639_), .A3(new_n555_), .A4(new_n875_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT126), .B1(new_n919_), .B2(new_n913_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n918_), .A2(new_n920_), .A3(new_n904_), .A4(new_n905_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n921_), .ZN(G1354gat));
  INV_X1    g721(.A(new_n898_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(KEYINPUT127), .A3(new_n647_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n898_), .B2(new_n674_), .ZN(new_n926_));
  INV_X1    g725(.A(G218gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n924_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n923_), .A2(G218gat), .A3(new_n681_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1355gat));
endmodule


