//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(G228gat), .ZN(new_n202_));
  INV_X1    g001(.A(G233gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  NOR3_X1   g004(.A1(new_n205_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(G204gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT89), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT21), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT88), .B1(new_n205_), .B2(G197gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT88), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(new_n207_), .A3(G204gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n205_), .A2(G197gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n212_), .A2(new_n215_), .A3(new_n211_), .A4(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT89), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT87), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G197gat), .B(G204gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(new_n211_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n205_), .A2(G197gat), .ZN(new_n223_));
  OAI211_X1 g022(.A(KEYINPUT87), .B(KEYINPUT21), .C1(new_n223_), .C2(new_n208_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT90), .ZN(new_n225_));
  INV_X1    g024(.A(G218gat), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n226_), .A2(G211gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(G211gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n225_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G211gat), .B(G218gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT90), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n222_), .A2(new_n224_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n231_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n211_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n219_), .A2(new_n232_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT84), .ZN(new_n238_));
  AND2_X1   g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G155gat), .ZN(new_n242_));
  INV_X1    g041(.A(G162gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT84), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT83), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n251_), .A2(G141gat), .A3(G148gat), .ZN(new_n252_));
  INV_X1    g051(.A(G141gat), .ZN(new_n253_));
  INV_X1    g052(.A(G148gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT3), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n250_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n247_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n245_), .A2(KEYINPUT1), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(G155gat), .A3(G162gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n262_), .A3(new_n244_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n253_), .A2(new_n254_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n237_), .B1(new_n259_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n204_), .B1(new_n236_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT91), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT91), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n270_), .B(new_n204_), .C1(new_n236_), .C2(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n234_), .A2(new_n235_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n217_), .B(new_n210_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n222_), .A2(new_n224_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n233_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n273_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT3), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n251_), .B1(G141gat), .B2(G148gat), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n278_), .A2(new_n279_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n280_));
  AND3_X1   g079(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n264_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n283_), .B2(KEYINPUT83), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n280_), .A2(new_n284_), .B1(new_n241_), .B2(new_n246_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT85), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT85), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n259_), .A2(new_n288_), .A3(new_n266_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  OAI221_X1 g089(.A(new_n277_), .B1(new_n202_), .B2(new_n203_), .C1(new_n290_), .C2(new_n237_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n272_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G78gat), .B(G106gat), .Z(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n272_), .A2(new_n291_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n290_), .A2(new_n237_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G22gat), .B(G50gat), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n299_), .B1(new_n290_), .B2(new_n237_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n301_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT92), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n303_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT92), .B1(new_n310_), .B2(new_n305_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n297_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n310_), .A2(KEYINPUT92), .A3(new_n305_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G8gat), .B(G36gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT18), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT24), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT94), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  INV_X1    g123(.A(G176gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT94), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n321_), .A2(new_n327_), .A3(KEYINPUT24), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G183gat), .ZN(new_n330_));
  INV_X1    g129(.A(G190gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT23), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(G183gat), .A3(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n326_), .A2(KEYINPUT24), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT25), .B(G183gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n329_), .A2(new_n335_), .A3(new_n336_), .A4(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n333_), .B1(G183gat), .B2(G190gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n334_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n333_), .A2(KEYINPUT78), .A3(G183gat), .A4(G190gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n321_), .A2(KEYINPUT77), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(G169gat), .A3(G176gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n324_), .A2(KEYINPUT22), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n324_), .A2(KEYINPUT22), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n350_), .B1(new_n354_), .B2(new_n325_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n340_), .B1(new_n346_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT20), .B1(new_n277_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n343_), .A2(new_n344_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n332_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n336_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n336_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT79), .B1(new_n345_), .B2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n347_), .A2(new_n349_), .A3(new_n326_), .A4(KEYINPUT24), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n339_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n330_), .A2(new_n331_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n350_), .B1(new_n335_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT80), .B1(new_n352_), .B2(new_n353_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372_));
  AOI21_X1  g171(.A(G176gat), .B1(new_n351_), .B2(new_n372_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n370_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n369_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n219_), .A2(new_n232_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n367_), .A2(new_n376_), .B1(new_n377_), .B2(new_n273_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n379_), .B(KEYINPUT19), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n358_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n380_), .B(KEYINPUT93), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT20), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n277_), .B2(new_n357_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n236_), .A2(new_n367_), .A3(new_n376_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n384_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n320_), .B1(new_n382_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n367_), .A2(new_n376_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(new_n277_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n360_), .A2(new_n368_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n339_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n392_), .A2(new_n355_), .B1(new_n393_), .B2(new_n329_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT20), .B1(new_n236_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n383_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n277_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n385_), .B1(new_n236_), .B2(new_n394_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n398_), .A3(new_n380_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(new_n399_), .A3(new_n319_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n389_), .A2(KEYINPUT95), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT95), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n403_), .B(new_n320_), .C1(new_n382_), .C2(new_n388_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n391_), .A2(new_n395_), .A3(new_n383_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n380_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n320_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(KEYINPUT27), .A3(new_n400_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n315_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G227gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(G15gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT30), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n390_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n418_));
  XOR2_X1   g217(.A(G127gat), .B(G134gat), .Z(new_n419_));
  XOR2_X1   g218(.A(G113gat), .B(G120gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT31), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n418_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(new_n422_), .B2(new_n421_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n417_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G43gat), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n427_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G1gat), .B(G29gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(G85gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT0), .B(G57gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n432_), .B(new_n433_), .Z(new_n434_));
  XOR2_X1   g233(.A(new_n419_), .B(new_n420_), .Z(new_n435_));
  NAND3_X1  g234(.A1(new_n287_), .A2(new_n289_), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n421_), .A2(new_n259_), .A3(new_n266_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(KEYINPUT4), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n287_), .A2(new_n289_), .A3(new_n441_), .A4(new_n435_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n436_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n434_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n434_), .A3(new_n444_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n430_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n412_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n401_), .A2(new_n404_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n447_), .A2(KEYINPUT33), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n443_), .A2(new_n454_), .A3(new_n434_), .A4(new_n444_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n436_), .A2(KEYINPUT4), .A3(new_n437_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n442_), .A2(new_n439_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n436_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n434_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT96), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT96), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n460_), .A4(new_n459_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n453_), .A2(new_n455_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n452_), .A2(new_n466_), .A3(KEYINPUT97), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT97), .B1(new_n452_), .B2(new_n466_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT32), .B(new_n319_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n319_), .A2(KEYINPUT32), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n396_), .A2(new_n399_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n447_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n469_), .B(new_n471_), .C1(new_n472_), .C2(new_n445_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n467_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT98), .B1(new_n475_), .B2(new_n315_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n452_), .A2(new_n466_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT97), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n474_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n452_), .A2(new_n466_), .A3(KEYINPUT97), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n315_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT98), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n312_), .A2(new_n314_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(new_n448_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n410_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n476_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n451_), .B1(new_n488_), .B2(new_n430_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G29gat), .B(G36gat), .Z(new_n490_));
  XOR2_X1   g289(.A(G43gat), .B(G50gat), .Z(new_n491_));
  XOR2_X1   g290(.A(new_n490_), .B(new_n491_), .Z(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT15), .Z(new_n493_));
  XOR2_X1   g292(.A(KEYINPUT71), .B(G8gat), .Z(new_n494_));
  INV_X1    g293(.A(G1gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G1gat), .B(G8gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n493_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n502_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n492_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT75), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n492_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n507_), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n512_), .B(KEYINPUT73), .Z(new_n513_));
  INV_X1    g312(.A(new_n508_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n513_), .A2(KEYINPUT74), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT74), .B1(new_n513_), .B2(new_n514_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n510_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G169gat), .B(G197gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n510_), .B(new_n520_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT76), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n522_), .A2(new_n526_), .A3(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n505_), .B(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G71gat), .B(G78gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G57gat), .B(G64gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n531_), .B1(KEYINPUT11), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT67), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(KEYINPUT11), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n530_), .B(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G127gat), .B(G155gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT16), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G183gat), .B(G211gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(KEYINPUT72), .A2(KEYINPUT17), .ZN(new_n542_));
  OR3_X1    g341(.A1(new_n537_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  MUX2_X1   g342(.A(new_n542_), .B(KEYINPUT17), .S(new_n541_), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n537_), .A2(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT8), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT6), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT66), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT7), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n553_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G85gat), .B(G92gat), .Z(new_n559_));
  AOI21_X1  g358(.A(new_n550_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n550_), .A2(KEYINPUT65), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n550_), .A2(KEYINPUT65), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n559_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT10), .B(G99gat), .Z(new_n571_));
  INV_X1    g370(.A(G106gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n569_), .A2(new_n570_), .A3(new_n552_), .A4(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n565_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT35), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n575_), .A2(new_n506_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n565_), .A2(new_n574_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n493_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n580_), .B(new_n582_), .C1(new_n576_), .C2(new_n579_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  OAI22_X1  g383(.A1(new_n581_), .A2(new_n492_), .B1(KEYINPUT35), .B2(new_n578_), .ZN(new_n585_));
  OAI211_X1 g384(.A(KEYINPUT35), .B(new_n578_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT69), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n588_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n583_), .A2(new_n586_), .A3(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n589_), .B1(new_n588_), .B2(new_n593_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n549_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n588_), .A2(new_n593_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT36), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n600_), .A2(new_n595_), .A3(new_n594_), .A4(new_n548_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n547_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n581_), .A2(new_n536_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n581_), .A2(new_n536_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(KEYINPUT12), .A3(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(KEYINPUT12), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(G230gat), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n203_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT5), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n612_), .A2(new_n614_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n610_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n618_), .B1(new_n621_), .B2(new_n613_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT68), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(KEYINPUT13), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n626_));
  NAND3_X1  g425(.A1(new_n620_), .A2(new_n622_), .A3(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NOR4_X1   g427(.A1(new_n489_), .A2(new_n528_), .A3(new_n603_), .A4(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n495_), .A3(new_n448_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n630_), .A2(new_n631_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n634_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n600_), .A2(KEYINPUT99), .A3(new_n595_), .A4(new_n594_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n489_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n625_), .A2(new_n627_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n524_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(new_n547_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n495_), .B1(new_n643_), .B2(new_n448_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n632_), .A2(new_n633_), .A3(new_n644_), .ZN(G1324gat));
  NAND3_X1  g444(.A1(new_n629_), .A2(new_n410_), .A3(new_n494_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n643_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G8gat), .B1(new_n647_), .B2(new_n486_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(KEYINPUT39), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(KEYINPUT39), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT40), .B(new_n646_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  INV_X1    g454(.A(new_n430_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n414_), .B1(new_n643_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n629_), .A2(new_n414_), .A3(new_n656_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT100), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n658_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n661_), .A3(new_n662_), .ZN(G1326gat));
  NOR2_X1   g462(.A1(new_n484_), .A2(G22gat), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT103), .Z(new_n665_));
  NAND2_X1  g464(.A1(new_n629_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n643_), .A2(new_n315_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G22gat), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT102), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(KEYINPUT102), .ZN(new_n670_));
  XOR2_X1   g469(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n666_), .B1(new_n672_), .B2(new_n673_), .ZN(G1327gat));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675_));
  NAND2_X1  g474(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n598_), .A2(new_n601_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n489_), .B2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n487_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n475_), .A2(KEYINPUT98), .A3(new_n315_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n430_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n451_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n681_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n676_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n682_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n641_), .A2(new_n546_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n690_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT44), .B1(new_n690_), .B2(new_n691_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n448_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G29gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n489_), .A2(new_n528_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n638_), .A2(new_n547_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n628_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n448_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n700_), .A2(G29gat), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n675_), .B1(new_n696_), .B2(new_n703_), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT105), .B(new_n702_), .C1(new_n695_), .C2(G29gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(new_n700_), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n410_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n692_), .A2(new_n693_), .A3(new_n486_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n712_), .B(KEYINPUT46), .C1(new_n708_), .C2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n713_), .A2(new_n708_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(new_n711_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(G1329gat));
  AOI21_X1  g517(.A(G43gat), .B1(new_n707_), .B2(new_n656_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n656_), .A2(G43gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n694_), .B2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT47), .Z(G1330gat));
  OR3_X1    g521(.A1(new_n700_), .A2(G50gat), .A3(new_n484_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n679_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n681_), .B(new_n677_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n691_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n690_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n728_), .A2(KEYINPUT107), .A3(new_n315_), .A4(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(G50gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n315_), .A3(new_n729_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT108), .B1(new_n731_), .B2(new_n734_), .ZN(new_n735_));
  AND4_X1   g534(.A1(KEYINPUT108), .A2(new_n734_), .A3(G50gat), .A4(new_n730_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n723_), .B1(new_n735_), .B2(new_n736_), .ZN(G1331gat));
  NOR2_X1   g536(.A1(new_n489_), .A2(new_n524_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n603_), .A2(new_n640_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n701_), .B1(new_n740_), .B2(KEYINPUT109), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(KEYINPUT109), .B2(new_n740_), .ZN(new_n742_));
  INV_X1    g541(.A(G57gat), .ZN(new_n743_));
  AND4_X1   g542(.A1(new_n528_), .A2(new_n639_), .A3(new_n628_), .A4(new_n546_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n701_), .A2(new_n743_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n742_), .A2(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(G64gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n744_), .B2(new_n410_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT48), .Z(new_n749_));
  INV_X1    g548(.A(new_n740_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n747_), .A3(new_n410_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n744_), .B2(new_n656_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT49), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n750_), .A2(new_n753_), .A3(new_n656_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1334gat));
  INV_X1    g556(.A(G78gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n744_), .B2(new_n315_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n750_), .A2(new_n758_), .A3(new_n315_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1335gat));
  NOR4_X1   g562(.A1(new_n489_), .A2(new_n698_), .A3(new_n524_), .A4(new_n640_), .ZN(new_n764_));
  INV_X1    g563(.A(G85gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n448_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n524_), .A2(new_n546_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n628_), .B2(new_n768_), .ZN(new_n769_));
  AND4_X1   g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n627_), .A4(new_n625_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n690_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n690_), .A2(KEYINPUT112), .A3(new_n772_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n701_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n766_), .B1(new_n777_), .B2(new_n765_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1336gat));
  INV_X1    g579(.A(G92gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n764_), .A2(new_n781_), .A3(new_n410_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n486_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n781_), .ZN(G1337gat));
  NAND3_X1  g583(.A1(new_n764_), .A2(new_n656_), .A3(new_n571_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n430_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n786_));
  INV_X1    g585(.A(G99gat), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT115), .B(new_n785_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790_));
  INV_X1    g589(.A(new_n785_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT112), .B1(new_n690_), .B2(new_n772_), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n774_), .B(new_n771_), .C1(new_n682_), .C2(new_n689_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n656_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n791_), .B1(new_n794_), .B2(G99gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n790_), .B1(new_n795_), .B2(KEYINPUT115), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n795_), .B2(new_n790_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n789_), .B1(new_n796_), .B2(new_n798_), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n764_), .A2(new_n572_), .A3(new_n315_), .ZN(new_n800_));
  OAI21_X1  g599(.A(G106gat), .B1(new_n773_), .B2(new_n484_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n801_), .A2(KEYINPUT52), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(KEYINPUT52), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n800_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n800_), .B(new_n805_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1339gat));
  NOR3_X1   g608(.A1(new_n412_), .A2(new_n701_), .A3(new_n430_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n524_), .A2(new_n620_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n608_), .A2(new_n611_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n621_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n619_), .B1(new_n621_), .B2(new_n814_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n812_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n621_), .A2(new_n814_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n611_), .B2(new_n608_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n816_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n811_), .B1(new_n818_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n513_), .A2(new_n509_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n509_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n520_), .B1(new_n504_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n523_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n622_), .B2(new_n620_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n637_), .B1(new_n822_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  INV_X1    g629(.A(new_n620_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n815_), .A2(new_n817_), .A3(new_n812_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n816_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n681_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n818_), .A2(new_n821_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT58), .A3(new_n832_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n829_), .A2(new_n830_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT57), .B(new_n637_), .C1(new_n822_), .C2(new_n828_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n546_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n602_), .A2(new_n528_), .A3(new_n640_), .A4(new_n843_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n602_), .A2(new_n528_), .A3(new_n640_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT59), .B(new_n810_), .C1(new_n842_), .C2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n835_), .A2(new_n836_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n688_), .A3(new_n839_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n831_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n828_), .B1(new_n838_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n830_), .B1(new_n854_), .B2(new_n638_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n855_), .A3(new_n841_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n848_), .B1(new_n856_), .B2(new_n547_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n810_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n850_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n528_), .B1(new_n849_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(G113gat), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n857_), .A2(new_n858_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n524_), .A2(new_n861_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT118), .B1(new_n862_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868_));
  OAI221_X1 g667(.A(new_n868_), .B1(new_n864_), .B2(new_n865_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1340gat));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n640_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n863_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n871_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n640_), .B1(new_n849_), .B2(new_n859_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n871_), .ZN(G1341gat));
  INV_X1    g674(.A(G127gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n863_), .A2(new_n876_), .A3(new_n546_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n547_), .B1(new_n849_), .B2(new_n859_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n876_), .ZN(G1342gat));
  INV_X1    g678(.A(G134gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n863_), .A2(new_n880_), .A3(new_n638_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n681_), .B1(new_n849_), .B2(new_n859_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n880_), .ZN(G1343gat));
  INV_X1    g682(.A(new_n857_), .ZN(new_n884_));
  NOR4_X1   g683(.A1(new_n656_), .A2(new_n484_), .A3(new_n701_), .A4(new_n410_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n524_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n886_), .A2(new_n640_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n254_), .ZN(G1345gat));
  NOR2_X1   g690(.A1(new_n886_), .A2(new_n547_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT61), .B(G155gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n886_), .B2(new_n681_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n638_), .A2(new_n243_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n886_), .B2(new_n896_), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n857_), .A2(new_n486_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n450_), .A2(new_n315_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n524_), .A2(new_n354_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT119), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n898_), .A2(new_n524_), .A3(new_n899_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n904_), .A2(new_n905_), .A3(G169gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n904_), .B2(G169gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n903_), .B1(new_n906_), .B2(new_n907_), .ZN(G1348gat));
  NAND2_X1  g707(.A1(new_n900_), .A2(new_n628_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT120), .B(G176gat), .Z(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1349gat));
  AOI21_X1  g710(.A(G183gat), .B1(new_n900_), .B2(new_n546_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n337_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n898_), .A2(new_n913_), .A3(new_n546_), .A4(new_n899_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n914_), .A2(KEYINPUT121), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(KEYINPUT121), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n912_), .A2(new_n915_), .A3(new_n916_), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n900_), .A2(new_n338_), .A3(new_n638_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n900_), .A2(new_n688_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n331_), .ZN(G1351gat));
  INV_X1    g719(.A(new_n898_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n485_), .A2(new_n430_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n524_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT122), .B(G197gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1352gat));
  NAND2_X1  g725(.A1(new_n923_), .A2(new_n628_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g727(.A(new_n547_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT123), .Z(new_n930_));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n931_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n923_), .A2(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n931_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT125), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n934_), .B(new_n936_), .ZN(G1354gat));
  NOR4_X1   g736(.A1(new_n857_), .A2(new_n486_), .A3(new_n637_), .A4(new_n922_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  OR2_X1    g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G218gat), .B1(new_n938_), .B2(new_n939_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n681_), .A2(new_n226_), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n940_), .A2(new_n941_), .B1(new_n923_), .B2(new_n942_), .ZN(G1355gat));
endmodule


