//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT10), .B(G99gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT65), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(new_n211_), .B2(G106gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n216_), .A2(new_n217_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n213_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n213_), .A2(new_n215_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n216_), .A2(new_n217_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(KEYINPUT67), .A3(new_n213_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n212_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n209_), .ZN(new_n229_));
  INV_X1    g028(.A(G99gat), .ZN(new_n230_));
  INV_X1    g029(.A(G106gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT68), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT7), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n234_), .A2(new_n230_), .A3(new_n231_), .A4(KEYINPUT68), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n223_), .B1(new_n229_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT8), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(KEYINPUT69), .A3(new_n235_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT69), .B1(new_n233_), .B2(new_n235_), .ZN(new_n242_));
  NOR3_X1   g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n229_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n223_), .A2(KEYINPUT8), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n239_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n207_), .B1(new_n228_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT74), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n210_), .B(KEYINPUT65), .Z(new_n248_));
  AOI21_X1  g047(.A(new_n229_), .B1(new_n248_), .B2(new_n231_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT67), .B1(new_n226_), .B2(new_n213_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n213_), .ZN(new_n251_));
  AOI211_X1 g050(.A(new_n221_), .B(new_n251_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n249_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n242_), .A2(new_n229_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n240_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n244_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n255_), .A2(new_n256_), .B1(new_n238_), .B2(new_n237_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT74), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n207_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n228_), .A2(new_n245_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n247_), .A2(new_n260_), .B1(new_n261_), .B2(new_n206_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT34), .Z(new_n264_));
  XOR2_X1   g063(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT75), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n247_), .B2(new_n260_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n264_), .A2(new_n265_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n262_), .B(new_n266_), .C1(new_n268_), .C2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n259_), .B1(new_n258_), .B2(new_n207_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT15), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n206_), .B(new_n273_), .ZN(new_n274_));
  AOI211_X1 g073(.A(KEYINPUT74), .B(new_n274_), .C1(new_n253_), .C2(new_n257_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT75), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n261_), .A2(new_n206_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n278_), .A3(new_n269_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G190gat), .B(G218gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(G134gat), .B(G162gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT76), .B(KEYINPUT77), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(KEYINPUT36), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n271_), .A2(new_n279_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(KEYINPUT36), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n271_), .A2(new_n279_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT37), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n271_), .A2(new_n279_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n271_), .A2(new_n279_), .A3(new_n285_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT37), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G127gat), .B(G155gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT16), .ZN(new_n299_));
  XOR2_X1   g098(.A(G183gat), .B(G211gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT17), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT78), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G15gat), .B(G22gat), .ZN(new_n305_));
  INV_X1    g104(.A(G1gat), .ZN(new_n306_));
  INV_X1    g105(.A(G8gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT14), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G1gat), .B(G8gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G64gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G71gat), .B(G78gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(KEYINPUT11), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(KEYINPUT11), .ZN(new_n317_));
  INV_X1    g116(.A(new_n315_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n314_), .A2(KEYINPUT11), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n316_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT70), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n323_), .B(new_n316_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n313_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n321_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n313_), .A2(new_n328_), .ZN(new_n329_));
  AOI211_X1 g128(.A(new_n302_), .B(new_n301_), .C1(new_n313_), .C2(new_n328_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n304_), .A2(new_n327_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n297_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT79), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT20), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n338_));
  INV_X1    g137(.A(G169gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT22), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT22), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(G176gat), .ZN(new_n343_));
  AND4_X1   g142(.A1(new_n338_), .A2(new_n340_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT22), .B(G169gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT84), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n353_));
  AND2_X1   g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n351_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(KEYINPUT23), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT24), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n350_), .A2(KEYINPUT24), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n365_), .B2(new_n362_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT25), .B(G183gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n369_));
  INV_X1    g168(.A(G190gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(KEYINPUT26), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT26), .B(G190gat), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n368_), .B(new_n371_), .C1(new_n372_), .C2(new_n369_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n349_), .A2(new_n358_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G218gat), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n375_), .A2(G211gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(G211gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT94), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G211gat), .B(G218gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G204gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT93), .B1(new_n382_), .B2(G197gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT93), .ZN(new_n384_));
  INV_X1    g183(.A(G197gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(G204gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(G197gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n378_), .A2(new_n381_), .A3(KEYINPUT21), .A4(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n382_), .A2(G197gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n385_), .A2(G204gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT21), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n392_), .B(new_n379_), .C1(new_n388_), .C2(KEYINPUT21), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n337_), .B1(new_n374_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n366_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n372_), .A2(new_n368_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n355_), .A3(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n399_));
  NAND2_X1  g198(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n354_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT96), .B(new_n357_), .C1(new_n401_), .C2(new_n360_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n351_), .B1(new_n346_), .B2(new_n343_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n405_));
  NOR2_X1   g204(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n359_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(KEYINPUT23), .B2(new_n359_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT96), .B1(new_n408_), .B2(new_n357_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n398_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n389_), .A2(new_n393_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n336_), .B1(new_n395_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT97), .ZN(new_n414_));
  INV_X1    g213(.A(new_n336_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT96), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n361_), .B2(new_n356_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n394_), .B1(new_n418_), .B2(new_n398_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n354_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n352_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n357_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n338_), .B1(new_n346_), .B2(new_n343_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n422_), .B(new_n350_), .C1(new_n423_), .C2(new_n344_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n396_), .A2(new_n373_), .A3(new_n408_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT20), .B1(new_n426_), .B2(new_n411_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n415_), .B1(new_n419_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT97), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G64gat), .B(G92gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT100), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT99), .B(KEYINPUT18), .Z(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n434_), .B(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT98), .B1(new_n410_), .B2(new_n411_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n337_), .B1(new_n426_), .B2(new_n411_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT98), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n418_), .A2(new_n394_), .A3(new_n440_), .A4(new_n398_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n438_), .A2(new_n439_), .A3(new_n336_), .A4(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n414_), .A2(new_n430_), .A3(new_n437_), .A4(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n395_), .A2(new_n336_), .A3(new_n412_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n418_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n439_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n446_), .B2(new_n336_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n437_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n443_), .A2(KEYINPUT27), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n442_), .B1(new_n413_), .B2(KEYINPUT97), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n428_), .A2(new_n429_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n448_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n443_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT27), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT103), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT103), .ZN(new_n457_));
  AOI211_X1 g256(.A(new_n457_), .B(KEYINPUT27), .C1(new_n453_), .C2(new_n443_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n450_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n424_), .A2(new_n425_), .A3(KEYINPUT30), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(G15gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G71gat), .ZN(new_n464_));
  INV_X1    g263(.A(G15gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n462_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G71gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(new_n230_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT30), .B1(new_n424_), .B2(new_n425_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n461_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n469_), .B(G99gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n460_), .B2(new_n471_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT85), .B(G43gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT31), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n479_), .A2(new_n480_), .A3(KEYINPUT88), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT88), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n473_), .A2(new_n475_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n477_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n482_), .B1(new_n485_), .B2(new_n478_), .ZN(new_n486_));
  INV_X1    g285(.A(G120gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G113gat), .ZN(new_n488_));
  INV_X1    g287(.A(G113gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G120gat), .ZN(new_n490_));
  INV_X1    g289(.A(G127gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(G134gat), .ZN(new_n492_));
  INV_X1    g291(.A(G134gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(G127gat), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n488_), .B(new_n490_), .C1(new_n492_), .C2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n490_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G127gat), .B(G134gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n502_));
  OAI22_X1  g301(.A1(new_n481_), .A2(new_n486_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT88), .B1(new_n479_), .B2(new_n480_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n485_), .A2(new_n482_), .A3(new_n478_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n501_), .A2(new_n502_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G1gat), .B(G29gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(G85gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT0), .B(G57gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(KEYINPUT102), .ZN(new_n513_));
  XOR2_X1   g312(.A(G155gat), .B(G162gat), .Z(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G141gat), .A2(G148gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT2), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G141gat), .A2(G148gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT3), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(KEYINPUT91), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n517_), .A2(new_n520_), .A3(new_n523_), .A4(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT92), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n528_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n514_), .B1(new_n525_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n521_), .A2(KEYINPUT89), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT89), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(G141gat), .B2(G148gat), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n532_), .A2(new_n518_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G155gat), .A2(G162gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G155gat), .A2(G162gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(KEYINPUT1), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT90), .B1(new_n536_), .B2(KEYINPUT1), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n536_), .A2(KEYINPUT90), .A3(KEYINPUT1), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n535_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n531_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544_));
  INV_X1    g343(.A(new_n502_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n500_), .A4(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT101), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT101), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n506_), .A2(new_n548_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n543_), .A2(new_n500_), .A3(new_n545_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n531_), .B(new_n542_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT4), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G225gat), .A2(G233gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n513_), .B1(new_n550_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n547_), .A2(new_n549_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n558_), .A2(KEYINPUT102), .A3(new_n553_), .A4(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n551_), .A2(new_n552_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n554_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n512_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n512_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n394_), .B1(KEYINPUT29), .B2(new_n543_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n543_), .A2(KEYINPUT29), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT28), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n568_), .A2(new_n569_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n567_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n567_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n543_), .A2(KEYINPUT29), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT28), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n576_), .A3(new_n570_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G228gat), .A2(G233gat), .ZN(new_n578_));
  INV_X1    g377(.A(G78gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n231_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G22gat), .B(G50gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n573_), .A2(new_n577_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n508_), .A2(new_n566_), .A3(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n459_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n512_), .B1(new_n561_), .B2(new_n555_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n553_), .A2(new_n554_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n589_), .B1(new_n550_), .B2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n453_), .A2(new_n443_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n564_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT33), .B1(new_n560_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n595_));
  AOI211_X1 g394(.A(new_n595_), .B(new_n564_), .C1(new_n557_), .C2(new_n559_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n592_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n437_), .A2(KEYINPUT32), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n414_), .A2(new_n598_), .A3(new_n442_), .A4(new_n430_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n447_), .A2(KEYINPUT32), .A3(new_n437_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n559_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n553_), .A2(new_n555_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT102), .B1(new_n603_), .B2(new_n558_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n562_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n512_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n593_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n601_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n586_), .B1(new_n597_), .B2(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n563_), .A2(new_n565_), .A3(new_n586_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n611_), .B(new_n450_), .C1(new_n456_), .C2(new_n458_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n508_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n588_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT64), .Z(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n253_), .A2(new_n257_), .A3(new_n325_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n325_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n618_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT5), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n328_), .A2(KEYINPUT12), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n228_), .B2(new_n245_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n619_), .B(new_n629_), .C1(new_n621_), .C2(KEYINPUT12), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n622_), .B(new_n626_), .C1(new_n630_), .C2(new_n618_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n626_), .B(KEYINPUT71), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n629_), .A2(new_n619_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT12), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n636_), .B1(new_n261_), .B2(new_n325_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n617_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n634_), .B1(new_n638_), .B2(new_n622_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT13), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(KEYINPUT72), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(KEYINPUT72), .ZN(new_n642_));
  OAI22_X1  g441(.A1(new_n632_), .A2(new_n639_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n622_), .B1(new_n630_), .B2(new_n618_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n633_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n642_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n631_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT80), .ZN(new_n649_));
  INV_X1    g448(.A(new_n311_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n206_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n311_), .A2(new_n205_), .A3(new_n204_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n649_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n207_), .A2(new_n311_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n654_), .A3(new_n651_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n657_), .A2(new_n649_), .A3(new_n654_), .A4(new_n651_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(KEYINPUT81), .A3(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(G113gat), .B(G141gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(G169gat), .B(G197gat), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n662_), .B(new_n663_), .Z(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n661_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n661_), .A2(new_n665_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n648_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n615_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n333_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n566_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n306_), .A3(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT105), .B1(new_n286_), .B2(new_n288_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n292_), .A2(new_n293_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n615_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n331_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n669_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G1gat), .B1(new_n683_), .B2(new_n566_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT106), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n675_), .A2(new_n685_), .ZN(G1324gat));
  NAND3_X1  g485(.A1(new_n671_), .A2(new_n307_), .A3(new_n459_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n680_), .A2(new_n459_), .A3(new_n682_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT39), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(G8gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n688_), .B2(G8gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n687_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1325gat));
  NAND3_X1  g494(.A1(new_n671_), .A2(new_n465_), .A3(new_n508_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n680_), .A2(new_n508_), .A3(new_n682_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT41), .B1(new_n697_), .B2(G15gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT108), .ZN(G1326gat));
  XOR2_X1   g501(.A(new_n586_), .B(KEYINPUT109), .Z(new_n703_));
  OAI21_X1  g502(.A(G22gat), .B1(new_n683_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT42), .ZN(new_n705_));
  INV_X1    g504(.A(G22gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n703_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n671_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1327gat));
  AND2_X1   g508(.A1(new_n676_), .A2(new_n678_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(new_n331_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n670_), .A2(new_n711_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n712_), .A2(G29gat), .A3(new_n566_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n648_), .A2(new_n681_), .A3(new_n668_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  XOR2_X1   g514(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n588_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n450_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n454_), .A2(new_n455_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n457_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n454_), .A2(KEYINPUT103), .A3(new_n455_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n601_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n608_), .A2(new_n595_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n565_), .A2(KEYINPUT33), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n728_), .B2(new_n592_), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n723_), .A2(new_n611_), .B1(new_n729_), .B2(new_n586_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n718_), .B1(new_n730_), .B2(new_n508_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n717_), .B1(new_n731_), .B2(new_n296_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n508_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n733_), .B(new_n296_), .C1(new_n734_), .C2(new_n588_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n715_), .B1(new_n732_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(KEYINPUT111), .A3(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n716_), .B1(new_n615_), .B2(new_n297_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n714_), .B1(new_n741_), .B2(new_n735_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n742_), .B2(KEYINPUT44), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n739_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n738_), .B(new_n714_), .C1(new_n741_), .C2(new_n735_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n566_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(G29gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n745_), .B1(new_n744_), .B2(new_n747_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n713_), .B1(new_n749_), .B2(new_n750_), .ZN(G1328gat));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(KEYINPUT46), .ZN(new_n753_));
  INV_X1    g552(.A(G36gat), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT44), .B(new_n715_), .C1(new_n732_), .C2(new_n736_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n459_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n754_), .B1(new_n744_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n459_), .A2(new_n754_), .ZN(new_n759_));
  OR3_X1    g558(.A1(new_n712_), .A2(KEYINPUT45), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT45), .B1(new_n712_), .B2(new_n759_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n753_), .B1(new_n758_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n753_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n756_), .B1(new_n743_), .B2(new_n739_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n765_), .B(new_n762_), .C1(new_n766_), .C2(new_n754_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(G1329gat));
  NAND2_X1  g567(.A1(new_n508_), .A2(G43gat), .ZN(new_n769_));
  AOI211_X1 g568(.A(new_n746_), .B(new_n769_), .C1(new_n739_), .C2(new_n743_), .ZN(new_n770_));
  INV_X1    g569(.A(G43gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n712_), .B2(new_n614_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT47), .B1(new_n770_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n744_), .A2(new_n755_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n775_), .B(new_n772_), .C1(new_n776_), .C2(new_n769_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(G1330gat));
  INV_X1    g577(.A(new_n712_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G50gat), .B1(new_n779_), .B2(new_n707_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n776_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n586_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(G50gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n780_), .B1(new_n781_), .B2(new_n783_), .ZN(G1331gat));
  INV_X1    g583(.A(new_n648_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n615_), .A2(new_n668_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n333_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(G57gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n672_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n668_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n680_), .A2(new_n331_), .A3(new_n785_), .A4(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G57gat), .B1(new_n791_), .B2(new_n566_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n792_), .ZN(G1332gat));
  OAI21_X1  g592(.A(G64gat), .B1(new_n791_), .B2(new_n723_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT48), .ZN(new_n795_));
  INV_X1    g594(.A(G64gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n796_), .A3(new_n459_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1333gat));
  OAI21_X1  g597(.A(G71gat), .B1(new_n791_), .B2(new_n614_), .ZN(new_n799_));
  XOR2_X1   g598(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n787_), .A2(new_n467_), .A3(new_n508_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1334gat));
  OAI21_X1  g602(.A(G78gat), .B1(new_n791_), .B2(new_n703_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT50), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n787_), .A2(new_n579_), .A3(new_n707_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(G1335gat));
  NOR3_X1   g606(.A1(new_n710_), .A2(new_n331_), .A3(new_n648_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n786_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G85gat), .B1(new_n810_), .B2(new_n672_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n785_), .A2(new_n681_), .A3(new_n790_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n741_), .B2(new_n735_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n672_), .A2(G85gat), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(KEYINPUT115), .Z(new_n815_));
  AOI21_X1  g614(.A(new_n811_), .B1(new_n813_), .B2(new_n815_), .ZN(G1336gat));
  INV_X1    g615(.A(G92gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n810_), .A2(new_n817_), .A3(new_n459_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n813_), .A2(new_n459_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n817_), .ZN(G1337gat));
  NOR2_X1   g619(.A1(new_n614_), .A2(new_n211_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT116), .B1(new_n810_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823_));
  INV_X1    g622(.A(new_n821_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n809_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT117), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n230_), .B1(new_n813_), .B2(new_n508_), .ZN(new_n827_));
  OR3_X1    g626(.A1(new_n826_), .A2(new_n827_), .A3(KEYINPUT51), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT51), .B1(new_n826_), .B2(new_n827_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1338gat));
  NAND3_X1  g629(.A1(new_n810_), .A2(new_n231_), .A3(new_n782_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n813_), .A2(new_n782_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(G106gat), .ZN(new_n834_));
  AOI211_X1 g633(.A(KEYINPUT52), .B(new_n231_), .C1(new_n813_), .C2(new_n782_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT53), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n831_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1339gat));
  XOR2_X1   g639(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n630_), .B2(new_n618_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n635_), .A2(KEYINPUT55), .A3(new_n637_), .A4(new_n617_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n630_), .A2(new_n618_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n633_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n633_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n632_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n645_), .A2(new_n631_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n665_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n657_), .A2(new_n651_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n655_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n651_), .A2(new_n654_), .A3(new_n652_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n664_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n854_), .A2(new_n858_), .ZN(new_n859_));
  AOI22_X1  g658(.A1(new_n851_), .A2(new_n852_), .B1(new_n853_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n841_), .B1(new_n860_), .B2(new_n679_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n850_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT56), .B1(new_n846_), .B2(new_n633_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n852_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n853_), .A2(new_n859_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n710_), .A2(new_n866_), .A3(KEYINPUT57), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n859_), .A2(new_n631_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n851_), .A2(KEYINPUT58), .A3(new_n868_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n296_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n861_), .A2(new_n867_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n681_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n331_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n643_), .B2(new_n647_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n289_), .A2(new_n877_), .A3(new_n295_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n289_), .A2(new_n877_), .A3(new_n295_), .A4(KEYINPUT118), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(KEYINPUT54), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n878_), .A2(new_n879_), .A3(new_n883_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n875_), .A2(new_n885_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n459_), .A2(new_n566_), .A3(new_n614_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n886_), .A2(new_n586_), .A3(new_n887_), .A4(new_n888_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n886_), .A2(new_n586_), .A3(new_n887_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(G113gat), .B1(new_n892_), .B2(new_n790_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n489_), .A3(new_n668_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1340gat));
  OAI21_X1  g694(.A(G120gat), .B1(new_n892_), .B2(new_n648_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n890_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n487_), .B1(new_n648_), .B2(KEYINPUT60), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(KEYINPUT60), .B2(new_n487_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n896_), .B1(new_n897_), .B2(new_n899_), .ZN(G1341gat));
  OAI21_X1  g699(.A(G127gat), .B1(new_n892_), .B2(new_n681_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n882_), .A2(new_n884_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n681_), .B2(new_n874_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n903_), .A2(new_n782_), .A3(new_n681_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n904_), .A2(new_n491_), .A3(new_n887_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n901_), .A2(new_n905_), .ZN(G1342gat));
  OAI21_X1  g705(.A(G134gat), .B1(new_n892_), .B2(new_n297_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n890_), .A2(new_n493_), .A3(new_n679_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1343gat));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n459_), .A2(new_n566_), .A3(new_n586_), .A4(new_n508_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n910_), .B1(new_n903_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n913_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n886_), .A2(KEYINPUT123), .A3(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n668_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n785_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n331_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT61), .B(G155gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1346gat));
  INV_X1    g723(.A(G162gat), .ZN(new_n925_));
  AOI211_X1 g724(.A(new_n925_), .B(new_n297_), .C1(new_n914_), .C2(new_n916_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n710_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n928_), .B2(G162gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(KEYINPUT123), .B1(new_n886_), .B2(new_n915_), .ZN(new_n930_));
  AOI211_X1 g729(.A(new_n910_), .B(new_n913_), .C1(new_n875_), .C2(new_n885_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n679_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n932_), .A2(KEYINPUT124), .A3(new_n925_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n926_), .B1(new_n929_), .B2(new_n933_), .ZN(G1347gat));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n508_), .A2(new_n566_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n707_), .A2(new_n723_), .A3(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n886_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n790_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n935_), .B1(new_n939_), .B2(new_n339_), .ZN(new_n940_));
  OAI211_X1 g739(.A(KEYINPUT62), .B(G169gat), .C1(new_n938_), .C2(new_n790_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n346_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n940_), .A2(new_n941_), .A3(new_n942_), .ZN(G1348gat));
  INV_X1    g742(.A(new_n938_), .ZN(new_n944_));
  AOI21_X1  g743(.A(G176gat), .B1(new_n944_), .B2(new_n785_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n903_), .A2(new_n782_), .ZN(new_n946_));
  NOR4_X1   g745(.A1(new_n723_), .A2(new_n648_), .A3(new_n936_), .A4(new_n343_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n945_), .B1(new_n946_), .B2(new_n947_), .ZN(G1349gat));
  NOR3_X1   g747(.A1(new_n938_), .A2(new_n368_), .A3(new_n681_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n904_), .A2(new_n566_), .A3(new_n459_), .A4(new_n508_), .ZN(new_n950_));
  INV_X1    g749(.A(G183gat), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n949_), .B1(new_n950_), .B2(new_n951_), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n938_), .B2(new_n297_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n679_), .A2(new_n372_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n938_), .B2(new_n954_), .ZN(G1351gat));
  NAND3_X1  g754(.A1(new_n459_), .A2(new_n611_), .A3(new_n614_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n903_), .A2(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n668_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n958_), .B1(KEYINPUT125), .B2(new_n385_), .ZN(new_n959_));
  XOR2_X1   g758(.A(KEYINPUT125), .B(G197gat), .Z(new_n960_));
  AOI21_X1  g759(.A(new_n959_), .B1(new_n958_), .B2(new_n960_), .ZN(G1352gat));
  NAND2_X1  g760(.A1(new_n957_), .A2(new_n785_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g762(.A(new_n681_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(KEYINPUT126), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n957_), .A2(new_n965_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(KEYINPUT127), .B2(new_n967_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n967_), .B(KEYINPUT127), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(new_n966_), .B2(new_n969_), .ZN(G1354gat));
  NAND3_X1  g769(.A1(new_n957_), .A2(new_n375_), .A3(new_n679_), .ZN(new_n971_));
  NOR3_X1   g770(.A1(new_n903_), .A2(new_n297_), .A3(new_n956_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n972_), .B2(new_n375_), .ZN(G1355gat));
endmodule


