//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_;
  XOR2_X1   g000(.A(G22gat), .B(G50gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OR2_X1    g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT83), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208_));
  INV_X1    g007(.A(G141gat), .ZN(new_n209_));
  INV_X1    g008(.A(G148gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n211_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT83), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n204_), .A2(new_n218_), .A3(new_n205_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n207_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n205_), .A2(KEYINPUT1), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G155gat), .A3(G162gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n223_), .A3(new_n204_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n209_), .A2(new_n210_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n212_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  OR3_X1    g026(.A1(new_n227_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT28), .B1(new_n227_), .B2(KEYINPUT29), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n229_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n203_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n233_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(new_n202_), .A3(new_n231_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT85), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G197gat), .B(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n239_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n238_), .A2(new_n239_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n238_), .A2(new_n239_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n241_), .B(new_n242_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n245_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n237_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G228gat), .ZN(new_n252_));
  INV_X1    g051(.A(G233gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n237_), .B(new_n250_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G78gat), .B(G106gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n234_), .B(new_n236_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n255_), .A2(new_n256_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n257_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT86), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n259_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT86), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n255_), .A2(KEYINPUT87), .A3(new_n256_), .A4(new_n258_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n265_), .A2(new_n267_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n234_), .A2(new_n236_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n262_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G225gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G127gat), .B(G134gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G113gat), .B(G120gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  XOR2_X1   g077(.A(KEYINPUT94), .B(KEYINPUT4), .Z(new_n279_));
  NAND3_X1  g078(.A1(new_n227_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n227_), .A2(new_n278_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n276_), .B(new_n277_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(new_n226_), .A3(new_n220_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n275_), .B(new_n280_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n281_), .A2(new_n283_), .A3(new_n274_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G1gat), .B(G29gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G57gat), .B(G85gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n281_), .A2(KEYINPUT4), .A3(new_n283_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n280_), .A2(new_n275_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n287_), .B(new_n295_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT27), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT89), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  INV_X1    g104(.A(new_n250_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT78), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT91), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(KEYINPUT24), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n313_), .B2(KEYINPUT24), .ZN(new_n317_));
  OR3_X1    g116(.A1(new_n312_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT92), .ZN(new_n319_));
  INV_X1    g118(.A(G183gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT25), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G183gat), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n321_), .A2(new_n323_), .A3(KEYINPUT90), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT90), .B1(new_n321_), .B2(new_n323_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G190gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n318_), .B(new_n319_), .C1(new_n326_), .C2(new_n328_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n324_), .A2(new_n328_), .A3(new_n325_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n312_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT92), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT23), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n329_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n313_), .A2(KEYINPUT79), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(G169gat), .A3(G176gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT81), .B(G176gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G169gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n334_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n306_), .B1(new_n338_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n312_), .A2(new_n335_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n327_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n350_), .A2(new_n334_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n312_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT24), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n353_), .A2(new_n354_), .A3(KEYINPUT80), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT80), .B1(new_n353_), .B2(new_n354_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n352_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n347_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n334_), .A2(KEYINPUT82), .A3(new_n346_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n345_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT20), .B1(new_n362_), .B2(new_n250_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n305_), .B1(new_n349_), .B2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G8gat), .B(G36gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n362_), .B2(new_n250_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n338_), .A2(new_n306_), .A3(new_n348_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n305_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n364_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n370_), .B1(new_n364_), .B2(new_n375_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n301_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n349_), .A2(new_n363_), .A3(new_n305_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n374_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n369_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n364_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(KEYINPUT27), .A3(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n273_), .A2(new_n300_), .A3(new_n378_), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n370_), .A2(KEYINPUT32), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n364_), .A2(new_n385_), .A3(new_n375_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n299_), .A2(new_n386_), .ZN(new_n387_));
  OR3_X1    g186(.A1(new_n349_), .A2(new_n363_), .A3(new_n305_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n380_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n385_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT33), .B1(new_n298_), .B2(KEYINPUT96), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT96), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n286_), .A2(new_n393_), .A3(new_n287_), .A4(new_n295_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n392_), .A2(KEYINPUT97), .A3(new_n394_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n286_), .A2(KEYINPUT33), .A3(new_n287_), .A4(new_n295_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n280_), .A2(new_n274_), .ZN(new_n401_));
  OAI221_X1 g200(.A(new_n293_), .B1(new_n284_), .B2(new_n274_), .C1(new_n296_), .C2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n376_), .A2(new_n377_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n391_), .B1(new_n399_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n384_), .B1(new_n405_), .B2(new_n273_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G43gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n362_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(new_n282_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(G15gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT30), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT31), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n410_), .B(new_n278_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n416_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n378_), .A2(new_n383_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT98), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT98), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n378_), .A2(new_n424_), .A3(new_n383_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n273_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n417_), .A2(new_n420_), .A3(new_n300_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n406_), .A2(new_n421_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT77), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n431_));
  XOR2_X1   g230(.A(KEYINPUT72), .B(G1gat), .Z(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT73), .B(G8gat), .Z(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G15gat), .B(G22gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(G1gat), .B(G8gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  OR3_X1    g236(.A1(new_n434_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G29gat), .B(G36gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G43gat), .B(G50gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n430_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n440_), .A2(KEYINPUT77), .A3(new_n444_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n444_), .B(KEYINPUT15), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n441_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n446_), .A2(new_n447_), .B1(new_n445_), .B2(new_n441_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n452_), .B1(new_n453_), .B2(new_n449_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G113gat), .B(G141gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G169gat), .B(G197gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n452_), .B(new_n457_), .C1(new_n453_), .C2(new_n449_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n429_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G85gat), .ZN(new_n463_));
  INV_X1    g262(.A(G92gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT9), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT9), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(G85gat), .A3(G92gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n470_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT65), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT65), .ZN(new_n480_));
  NOR4_X1   g279(.A1(new_n475_), .A2(new_n476_), .A3(new_n480_), .A4(G106gat), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n467_), .B(new_n474_), .C1(new_n479_), .C2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n483_));
  INV_X1    g282(.A(G99gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n478_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n470_), .A3(new_n473_), .A4(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT8), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n465_), .A2(new_n466_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n488_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT68), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n487_), .A2(new_n489_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT8), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n482_), .B1(new_n492_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT35), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G232gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT34), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n498_), .A2(new_n450_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT66), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n490_), .A2(new_n491_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n467_), .A2(new_n470_), .A3(new_n473_), .A4(new_n472_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n479_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n481_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n504_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n482_), .B(KEYINPUT66), .C1(new_n491_), .C2(new_n490_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n444_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n513_), .A2(KEYINPUT70), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(KEYINPUT70), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n503_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n502_), .A2(new_n499_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G190gat), .B(G218gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT71), .ZN(new_n520_));
  XOR2_X1   g319(.A(G134gat), .B(G162gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n513_), .B(KEYINPUT70), .ZN(new_n526_));
  INV_X1    g325(.A(new_n517_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n503_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n518_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n522_), .B(new_n523_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n518_), .B2(new_n528_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT37), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n518_), .A2(new_n528_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT37), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n518_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT74), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G71gat), .B(G78gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(new_n545_), .A3(KEYINPUT11), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n440_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n550_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n542_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n552_), .A2(new_n554_), .A3(new_n542_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT76), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G127gat), .B(G155gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G183gat), .B(G211gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n558_), .A2(KEYINPUT17), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n557_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n555_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n567_), .B2(KEYINPUT76), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n567_), .B2(new_n565_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n564_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n539_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT13), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT64), .Z(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n512_), .B2(new_n553_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n510_), .A2(new_n551_), .A3(new_n511_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n549_), .A2(KEYINPUT12), .A3(new_n550_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n498_), .A2(KEYINPUT69), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT69), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT68), .B1(new_n490_), .B2(new_n491_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n495_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n509_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n583_), .B1(new_n586_), .B2(new_n580_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n576_), .A2(new_n579_), .A3(new_n582_), .A4(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G120gat), .B(G148gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT5), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G176gat), .B(G204gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n577_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n512_), .A2(new_n553_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT67), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT67), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n512_), .A2(new_n597_), .A3(new_n553_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n594_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n575_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n588_), .B(new_n593_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT67), .B(new_n551_), .C1(new_n511_), .C2(new_n510_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n597_), .B1(new_n512_), .B2(new_n553_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n577_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n575_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n593_), .B1(new_n606_), .B2(new_n588_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n573_), .B1(new_n602_), .B2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n588_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n592_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(KEYINPUT13), .A3(new_n601_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n572_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n462_), .A2(new_n613_), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n614_), .A2(new_n432_), .A3(new_n300_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT99), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT99), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(KEYINPUT38), .A3(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n612_), .A2(new_n461_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n571_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n535_), .A2(new_n537_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n429_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(KEYINPUT101), .A3(new_n625_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n299_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G1gat), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n616_), .A2(new_n617_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(KEYINPUT102), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT102), .B1(new_n634_), .B2(new_n635_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n618_), .B(new_n633_), .C1(new_n636_), .C2(new_n637_), .ZN(G1324gat));
  INV_X1    g437(.A(new_n425_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n424_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n614_), .A2(new_n433_), .A3(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n622_), .A2(new_n641_), .A3(new_n625_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n644_), .A2(new_n645_), .A3(G8gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n644_), .B2(G8gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g448(.A(new_n421_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(G15gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT41), .B1(new_n650_), .B2(new_n413_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n614_), .A2(G15gat), .A3(new_n421_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT103), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n653_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n653_), .A2(new_n654_), .A3(KEYINPUT104), .A4(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1326gat));
  INV_X1    g460(.A(new_n273_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n614_), .A2(G22gat), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n273_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(G22gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n664_), .B2(G22gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(G1327gat));
  INV_X1    g467(.A(new_n571_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n619_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n539_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n421_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n376_), .A2(new_n377_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n403_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n673_), .A2(new_n397_), .A3(new_n674_), .A4(new_n398_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n387_), .A2(new_n390_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n662_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n672_), .B1(new_n678_), .B2(new_n384_), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n273_), .B(new_n427_), .C1(new_n423_), .C2(new_n425_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n671_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n273_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n273_), .A2(new_n300_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n422_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n421_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n662_), .B(new_n428_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n539_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n683_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n670_), .B1(new_n682_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT44), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(G29gat), .A3(new_n299_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n670_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT43), .B1(new_n681_), .B2(KEYINPUT105), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n689_), .A2(new_n690_), .A3(new_n683_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n624_), .A2(new_n669_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n612_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n462_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n300_), .ZN(new_n705_));
  OAI22_X1  g504(.A1(new_n694_), .A2(new_n701_), .B1(G29gat), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT106), .ZN(G1328gat));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n641_), .A2(KEYINPUT108), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n641_), .A2(KEYINPUT108), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n462_), .A2(new_n708_), .A3(new_n703_), .A4(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT45), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n642_), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n700_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT107), .B1(new_n715_), .B2(G36gat), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  AOI211_X1 g516(.A(new_n717_), .B(new_n708_), .C1(new_n714_), .C2(new_n700_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT46), .B(new_n713_), .C1(new_n716_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  XOR2_X1   g522(.A(KEYINPUT109), .B(G43gat), .Z(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n704_), .B2(new_n421_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n693_), .A2(G43gat), .A3(new_n672_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n701_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n693_), .A2(new_n273_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n701_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G50gat), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n701_), .A2(new_n730_), .A3(new_n729_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n662_), .A2(G50gat), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT111), .ZN(new_n735_));
  OAI22_X1  g534(.A1(new_n732_), .A2(new_n733_), .B1(new_n704_), .B2(new_n735_), .ZN(G1331gat));
  NAND2_X1  g535(.A1(new_n459_), .A2(new_n460_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n612_), .ZN(new_n738_));
  NOR4_X1   g537(.A1(new_n429_), .A2(new_n572_), .A3(new_n737_), .A4(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G57gat), .B1(new_n739_), .B2(new_n299_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n669_), .A2(new_n737_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n625_), .A2(new_n612_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G57gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n299_), .B2(KEYINPUT112), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(KEYINPUT112), .B2(new_n743_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n740_), .B1(new_n742_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(G64gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n739_), .A2(new_n747_), .A3(new_n711_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n742_), .A2(new_n711_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G64gat), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n753_));
  AND2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n752_), .A2(new_n753_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n748_), .B1(new_n754_), .B2(new_n755_), .ZN(G1333gat));
  INV_X1    g555(.A(G71gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n742_), .B2(new_n672_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT49), .Z(new_n759_));
  NAND3_X1  g558(.A1(new_n739_), .A2(new_n757_), .A3(new_n672_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1334gat));
  INV_X1    g560(.A(G78gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n742_), .B2(new_n273_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT50), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n739_), .A2(new_n762_), .A3(new_n273_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1335gat));
  NOR4_X1   g565(.A1(new_n429_), .A2(new_n737_), .A3(new_n738_), .A4(new_n702_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT115), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n463_), .A3(new_n299_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n682_), .A2(new_n691_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n738_), .A2(new_n737_), .A3(new_n571_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(new_n299_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n773_), .B2(new_n463_), .ZN(G1336gat));
  NAND3_X1  g573(.A1(new_n768_), .A2(new_n464_), .A3(new_n641_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n772_), .A2(new_n711_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n464_), .ZN(G1337gat));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n672_), .A3(new_n477_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n772_), .A2(new_n672_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n484_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g580(.A1(new_n770_), .A2(new_n273_), .A3(new_n771_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT116), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n770_), .A2(new_n784_), .A3(new_n273_), .A4(new_n771_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n478_), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n768_), .A2(new_n478_), .A3(new_n273_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n789_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n783_), .A2(new_n792_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n790_), .A2(new_n791_), .A3(new_n796_), .A4(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  NAND4_X1  g597(.A1(new_n608_), .A2(new_n611_), .A3(new_n461_), .A4(new_n571_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n799_), .A2(KEYINPUT118), .B1(new_n538_), .B2(new_n532_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n738_), .A2(new_n801_), .A3(new_n741_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n800_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n737_), .A2(new_n601_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n588_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n588_), .B2(new_n809_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n579_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(KEYINPUT55), .A4(new_n576_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT120), .B1(new_n588_), .B2(new_n809_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n579_), .A2(new_n595_), .A3(new_n582_), .A4(new_n587_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n575_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n592_), .B1(new_n812_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT56), .B(new_n592_), .C1(new_n812_), .C2(new_n819_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n807_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n449_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n448_), .A2(new_n825_), .A3(new_n451_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n826_), .B(new_n458_), .C1(new_n825_), .C2(new_n453_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n460_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n610_), .B2(new_n601_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n623_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n828_), .A2(new_n602_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n823_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n498_), .A2(new_n581_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n835_), .A2(new_n583_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(KEYINPUT55), .A3(new_n582_), .A4(new_n576_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n837_), .A2(KEYINPUT120), .B1(new_n575_), .B2(new_n817_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n815_), .C1(new_n811_), .C2(new_n810_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT56), .B1(new_n839_), .B2(new_n592_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n833_), .B1(new_n834_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(KEYINPUT58), .B(new_n833_), .C1(new_n834_), .C2(new_n840_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n671_), .A3(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT57), .B(new_n623_), .C1(new_n824_), .C2(new_n829_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n832_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n806_), .B1(new_n847_), .B2(new_n669_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n426_), .A2(new_n299_), .A3(new_n672_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(G113gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(new_n737_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n461_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n852_), .B1(new_n855_), .B2(new_n851_), .ZN(G1340gat));
  AOI21_X1  g655(.A(new_n738_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n857_));
  INV_X1    g656(.A(G120gat), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n738_), .A2(KEYINPUT60), .ZN(new_n859_));
  MUX2_X1   g658(.A(KEYINPUT60), .B(new_n859_), .S(new_n858_), .Z(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT121), .B1(new_n850_), .B2(new_n860_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n850_), .A2(KEYINPUT121), .A3(new_n860_), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n857_), .A2(new_n858_), .B1(new_n861_), .B2(new_n862_), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n850_), .A2(new_n864_), .A3(new_n571_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n669_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1342gat));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n850_), .A2(new_n868_), .A3(new_n624_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n539_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n868_), .ZN(G1343gat));
  NOR3_X1   g670(.A1(new_n672_), .A2(new_n662_), .A3(new_n300_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n709_), .A2(new_n710_), .A3(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT122), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n848_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n461_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n209_), .ZN(G1344gat));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n738_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n210_), .ZN(G1345gat));
  NOR2_X1   g678(.A1(new_n875_), .A2(new_n669_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT61), .B(G155gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n875_), .B2(new_n539_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n623_), .A2(G162gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n875_), .B2(new_n884_), .ZN(G1347gat));
  NAND3_X1  g684(.A1(new_n711_), .A2(new_n662_), .A3(new_n428_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n848_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888_), .B2(new_n461_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n887_), .A2(new_n737_), .A3(new_n344_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n890_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(G1348gat));
  NAND2_X1  g693(.A1(new_n887_), .A2(new_n612_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT123), .B1(new_n895_), .B2(new_n309_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n343_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n895_), .A2(KEYINPUT123), .A3(new_n309_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1349gat));
  NOR2_X1   g699(.A1(new_n888_), .A2(new_n669_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(G183gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n901_), .B2(new_n326_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n888_), .B2(new_n539_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n624_), .A2(new_n327_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT124), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n888_), .B2(new_n906_), .ZN(G1351gat));
  NAND4_X1  g706(.A1(new_n711_), .A2(new_n273_), .A3(new_n300_), .A4(new_n421_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n847_), .A2(new_n669_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n806_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n737_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n612_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g714(.A(new_n669_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n911_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT125), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n911_), .A2(new_n919_), .A3(new_n916_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  OR2_X1    g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1354gat));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n911_), .B2(new_n624_), .ZN(new_n925_));
  NOR4_X1   g724(.A1(new_n848_), .A2(KEYINPUT126), .A3(new_n623_), .A4(new_n908_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n925_), .A2(new_n926_), .A3(G218gat), .ZN(new_n927_));
  INV_X1    g726(.A(G218gat), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n539_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n911_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT127), .B1(new_n927_), .B2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n848_), .A2(new_n623_), .A3(new_n908_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n928_), .B1(new_n934_), .B2(new_n924_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n933_), .B(new_n930_), .C1(new_n935_), .C2(new_n926_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n932_), .A2(new_n936_), .ZN(G1355gat));
endmodule


