//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n204_), .B(new_n205_), .C1(new_n208_), .C2(KEYINPUT24), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(G169gat), .B2(G176gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT26), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT79), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n213_), .A2(KEYINPUT26), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(KEYINPUT79), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n204_), .B(new_n205_), .C1(G183gat), .C2(G190gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n206_), .A2(new_n207_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT22), .B(G169gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(new_n207_), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n212_), .A2(new_n219_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G227gat), .A2(G233gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G127gat), .ZN(new_n227_));
  INV_X1    g026(.A(G134gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G127gat), .A2(G134gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G113gat), .ZN(new_n232_));
  INV_X1    g031(.A(G120gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G113gat), .A2(G120gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n236_), .A3(KEYINPUT80), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n229_), .A2(new_n234_), .A3(new_n230_), .A4(new_n235_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT81), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n226_), .B(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT30), .B(G15gat), .Z(new_n246_));
  XNOR2_X1  g045(.A(G71gat), .B(G99gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT31), .B(G43gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n245_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n255_));
  INV_X1    g054(.A(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n256_), .ZN(new_n260_));
  INV_X1    g059(.A(G197gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n254_), .B1(new_n264_), .B2(KEYINPUT21), .ZN(new_n265_));
  AND2_X1   g064(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(G197gat), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(G204gat), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT21), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n268_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT89), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n268_), .A2(new_n271_), .A3(KEYINPUT89), .A4(new_n272_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT90), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n253_), .B(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n272_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(G190gat), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n217_), .A2(new_n283_), .B1(new_n211_), .B2(new_n208_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n209_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n284_), .A2(new_n285_), .B1(new_n223_), .B2(new_n220_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n224_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT20), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT19), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n277_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT20), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n292_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n224_), .B1(new_n281_), .B2(new_n277_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT93), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n224_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n282_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT93), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n299_), .A4(new_n301_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n293_), .A2(new_n298_), .A3(new_n304_), .A4(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT27), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT92), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n282_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n277_), .A2(KEYINPUT92), .A3(new_n281_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n287_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n306_), .A2(KEYINPUT20), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n292_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n224_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n286_), .B1(new_n277_), .B2(new_n281_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n300_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n292_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n298_), .B1(new_n316_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT101), .B1(new_n310_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n298_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n313_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT92), .B1(new_n277_), .B2(new_n281_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n286_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n303_), .A2(new_n300_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n320_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n290_), .A2(new_n292_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n324_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT101), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT27), .A4(new_n309_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n323_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n304_), .B(new_n308_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n324_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n309_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT102), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT102), .ZN(new_n340_));
  AOI211_X1 g139(.A(new_n340_), .B(KEYINPUT27), .C1(new_n336_), .C2(new_n309_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n334_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT82), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n344_), .A2(new_n346_), .B1(KEYINPUT83), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT83), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n343_), .A2(KEYINPUT82), .A3(new_n345_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n347_), .B2(KEYINPUT83), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .A4(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(KEYINPUT1), .B2(new_n355_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(KEYINPUT1), .B2(new_n355_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n344_), .A2(new_n352_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n354_), .A2(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  OR4_X1    g161(.A1(KEYINPUT98), .A2(new_n244_), .A3(KEYINPUT4), .A4(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT97), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT98), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n244_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT95), .B1(new_n244_), .B2(new_n362_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n354_), .A2(new_n358_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n360_), .A2(new_n361_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n371_), .A2(new_n243_), .A3(new_n372_), .A4(new_n241_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n237_), .A2(new_n242_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT96), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n362_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n367_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n363_), .B(new_n365_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT100), .B(G1gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n374_), .A2(new_n379_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n365_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n382_), .A2(new_n388_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n388_), .B1(new_n382_), .B2(new_n391_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n371_), .A2(KEYINPUT29), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n395_), .A2(KEYINPUT28), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(KEYINPUT28), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G22gat), .B(G50gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n396_), .A2(new_n397_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n404_));
  NAND2_X1  g203(.A1(new_n371_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n312_), .A2(new_n313_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G228gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT85), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G78gat), .B(G106gat), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n408_), .B(KEYINPUT86), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n371_), .A2(KEYINPUT84), .A3(KEYINPUT29), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT84), .B1(new_n371_), .B2(KEYINPUT29), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n282_), .B(new_n412_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n411_), .B1(new_n409_), .B2(new_n415_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n403_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n420_), .A2(new_n402_), .A3(new_n400_), .A4(new_n416_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n394_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n342_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n382_), .A2(new_n388_), .A3(new_n391_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n337_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n382_), .A2(KEYINPUT33), .A3(new_n388_), .A4(new_n391_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n388_), .B1(new_n389_), .B2(new_n365_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n363_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(new_n365_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n298_), .A2(KEYINPUT32), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n335_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n435_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n436_), .B(new_n437_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n422_), .B1(new_n433_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n252_), .B1(new_n424_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT103), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n342_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n334_), .B(KEYINPUT103), .C1(new_n339_), .C2(new_n341_), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n392_), .A2(new_n393_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(new_n422_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n442_), .A2(new_n251_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n440_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G120gat), .B(G148gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(new_n256_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT5), .B(G176gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G230gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT8), .ZN(new_n455_));
  XOR2_X1   g254(.A(G85gat), .B(G92gat), .Z(new_n456_));
  NOR2_X1   g255(.A1(G99gat), .A2(G106gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G99gat), .A2(G106gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n455_), .B(new_n456_), .C1(new_n459_), .C2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n456_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n459_), .B1(KEYINPUT65), .B2(new_n462_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n460_), .B(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n464_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n463_), .B1(new_n469_), .B2(new_n455_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G71gat), .B(G78gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(G57gat), .B(G64gat), .Z(new_n472_));
  INV_X1    g271(.A(KEYINPUT11), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G64gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n475_), .A2(new_n471_), .A3(KEYINPUT11), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G106gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(KEYINPUT10), .B(G99gat), .Z(new_n484_));
  AOI21_X1  g283(.A(new_n462_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n456_), .A2(KEYINPUT9), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G85gat), .A2(G92gat), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n485_), .B(new_n486_), .C1(KEYINPUT9), .C2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n470_), .A2(new_n482_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n462_), .A2(KEYINPUT65), .ZN(new_n490_));
  INV_X1    g289(.A(G99gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n483_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(new_n458_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n468_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n455_), .B1(new_n494_), .B2(new_n456_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n463_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n488_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n481_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n489_), .A2(new_n501_), .A3(KEYINPUT12), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT12), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n497_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n454_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n453_), .B1(new_n489_), .B2(new_n501_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n452_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n505_), .A2(new_n506_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n509_), .B2(new_n451_), .ZN(new_n510_));
  NOR4_X1   g309(.A1(new_n505_), .A2(KEYINPUT68), .A3(new_n506_), .A4(new_n452_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n507_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT13), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n502_), .A2(new_n504_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n453_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n506_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n516_), .A3(new_n451_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT68), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n509_), .A2(new_n508_), .A3(new_n451_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT13), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n507_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n513_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G29gat), .B(G36gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT15), .ZN(new_n527_));
  XOR2_X1   g326(.A(G29gat), .B(G36gat), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n525_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G43gat), .B(G50gat), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n524_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G1gat), .A2(G8gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT14), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n537_), .B1(new_n536_), .B2(KEYINPUT14), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n535_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G1gat), .B(G8gat), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n541_), .B(new_n535_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n527_), .A2(new_n534_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n544_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(new_n532_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT74), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n527_), .A2(new_n534_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n546_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT74), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n546_), .B(new_n532_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n553_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(KEYINPUT76), .B(new_n556_), .C1(new_n560_), .C2(new_n555_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT76), .ZN(new_n562_));
  INV_X1    g361(.A(new_n556_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n555_), .B1(new_n554_), .B2(new_n559_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G169gat), .B(G197gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT77), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n561_), .A2(new_n565_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT78), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n561_), .A2(new_n565_), .A3(new_n573_), .A4(new_n570_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n556_), .B(new_n569_), .C1(new_n560_), .C2(new_n555_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n523_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n447_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT36), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n470_), .A2(new_n488_), .A3(new_n526_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT69), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n590_));
  AOI211_X1 g389(.A(KEYINPUT70), .B(new_n590_), .C1(new_n497_), .C2(new_n549_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n587_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n584_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n594_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n582_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n596_), .A2(new_n592_), .A3(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT37), .B1(new_n595_), .B2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n593_), .A2(new_n597_), .A3(new_n582_), .A4(new_n594_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n583_), .B1(new_n596_), .B2(new_n592_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n546_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n500_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610_));
  INV_X1    g409(.A(G211gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT16), .B(G183gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n609_), .A2(KEYINPUT17), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT72), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n614_), .B(KEYINPUT17), .ZN(new_n617_));
  INV_X1    g416(.A(new_n609_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT73), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n619_), .B2(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n606_), .A2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n579_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n625_), .A2(G1gat), .A3(new_n394_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT105), .B1(new_n595_), .B2(new_n599_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n601_), .A2(new_n602_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n622_), .B(new_n632_), .C1(new_n440_), .C2(new_n446_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n513_), .A2(new_n522_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(KEYINPUT104), .A3(new_n576_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT104), .B1(new_n634_), .B2(new_n576_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n394_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n626_), .A2(new_n627_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n628_), .A2(new_n640_), .A3(new_n641_), .ZN(G1324gat));
  NAND2_X1  g441(.A1(new_n442_), .A2(new_n443_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n633_), .A2(new_n638_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n644_), .A2(new_n645_), .A3(G8gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n644_), .B2(G8gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n643_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(G8gat), .ZN(new_n649_));
  OAI22_X1  g448(.A1(new_n646_), .A2(new_n647_), .B1(new_n625_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g450(.A(G15gat), .B1(new_n639_), .B2(new_n252_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT41), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(KEYINPUT41), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n252_), .A2(G15gat), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n653_), .B(new_n654_), .C1(new_n625_), .C2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT106), .Z(G1326gat));
  INV_X1    g456(.A(new_n422_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G22gat), .B1(new_n639_), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n658_), .A2(G22gat), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n661_), .B(new_n662_), .C1(new_n625_), .C2(new_n663_), .ZN(G1327gat));
  INV_X1    g463(.A(new_n632_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n622_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n579_), .A2(new_n667_), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n668_), .A2(G29gat), .A3(new_n394_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n605_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n636_), .A2(new_n666_), .A3(new_n637_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT44), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n672_), .B1(new_n447_), .B2(new_n606_), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT43), .B(new_n605_), .C1(new_n440_), .C2(new_n446_), .ZN(new_n677_));
  OAI211_X1 g476(.A(KEYINPUT44), .B(new_n674_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n444_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n670_), .B(G29gat), .C1(new_n675_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n674_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n444_), .A3(new_n678_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n670_), .B1(new_n685_), .B2(G29gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n669_), .B1(new_n681_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT109), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n689_), .B(new_n669_), .C1(new_n681_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n684_), .A2(new_n643_), .A3(new_n678_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n648_), .A2(G36gat), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n694_), .A2(new_n447_), .A3(new_n667_), .A4(new_n578_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT45), .Z(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(KEYINPUT46), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT112), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n692_), .B2(G36gat), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT112), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n700_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n705_), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n678_), .A2(new_n643_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n684_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT111), .B(new_n707_), .C1(new_n710_), .C2(new_n696_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n706_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n703_), .A2(new_n712_), .ZN(G1329gat));
  NAND3_X1  g512(.A1(new_n678_), .A2(G43gat), .A3(new_n251_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n668_), .A2(new_n252_), .ZN(new_n715_));
  OAI22_X1  g514(.A1(new_n714_), .A2(new_n675_), .B1(G43gat), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g516(.A1(new_n678_), .A2(new_n422_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G50gat), .B1(new_n675_), .B2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n658_), .A2(G50gat), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT113), .Z(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n668_), .B2(new_n721_), .ZN(G1331gat));
  NAND2_X1  g521(.A1(new_n623_), .A2(new_n523_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n577_), .B1(new_n723_), .B2(KEYINPUT114), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(KEYINPUT114), .B2(new_n723_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n447_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n444_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n634_), .A2(new_n576_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n633_), .A2(G57gat), .A3(new_n444_), .A4(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(KEYINPUT115), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n730_), .A2(KEYINPUT115), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n728_), .A2(new_n731_), .A3(new_n732_), .ZN(G1332gat));
  NAND2_X1  g532(.A1(new_n633_), .A2(new_n729_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G64gat), .B1(new_n734_), .B2(new_n648_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT48), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n648_), .A2(G64gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n726_), .B2(new_n737_), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n734_), .B2(new_n252_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT49), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n252_), .A2(G71gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT116), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n726_), .B2(new_n742_), .ZN(G1334gat));
  OAI21_X1  g542(.A(G78gat), .B1(new_n734_), .B2(new_n658_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT50), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n658_), .A2(G78gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n726_), .B2(new_n746_), .ZN(G1335gat));
  NAND3_X1  g546(.A1(new_n447_), .A2(new_n667_), .A3(new_n729_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n444_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n676_), .A2(new_n677_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n729_), .A2(new_n622_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n444_), .A2(G85gat), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT117), .Z(new_n755_));
  AOI21_X1  g554(.A(new_n750_), .B1(new_n753_), .B2(new_n755_), .ZN(G1336gat));
  AOI21_X1  g555(.A(G92gat), .B1(new_n749_), .B2(new_n643_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n643_), .A2(G92gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n753_), .B2(new_n758_), .ZN(G1337gat));
  NAND2_X1  g558(.A1(new_n753_), .A2(new_n251_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G99gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n749_), .A2(new_n484_), .A3(new_n251_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n761_), .A2(new_n762_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n764_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(G1338gat));
  NAND3_X1  g566(.A1(new_n749_), .A2(new_n483_), .A3(new_n422_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n752_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(new_n422_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n483_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n768_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n768_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  NOR2_X1   g580(.A1(new_n643_), .A2(new_n252_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n444_), .A3(new_n658_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n548_), .A2(new_n552_), .A3(new_n558_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n569_), .B1(new_n557_), .B2(new_n553_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT121), .Z(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n575_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n520_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n514_), .A2(new_n453_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n515_), .A2(KEYINPUT55), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n505_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n790_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n451_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n505_), .A2(new_n792_), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT55), .B(new_n454_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n798_));
  OAI22_X1  g597(.A1(new_n797_), .A2(new_n798_), .B1(new_n453_), .B2(new_n514_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n452_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n789_), .B1(new_n796_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n605_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n802_), .B2(new_n801_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n795_), .B1(new_n794_), .B2(new_n451_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n452_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT120), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n799_), .A2(new_n808_), .A3(KEYINPUT56), .A4(new_n452_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n807_), .A2(new_n520_), .A3(new_n576_), .A4(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n512_), .A2(new_n788_), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT57), .B(new_n632_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n796_), .A2(new_n800_), .A3(new_n808_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n576_), .A2(new_n520_), .A3(new_n809_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n813_), .B1(new_n816_), .B2(new_n665_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n804_), .B1(new_n812_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT122), .B(new_n804_), .C1(new_n812_), .C2(new_n817_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n622_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n623_), .A2(new_n634_), .A3(new_n577_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT54), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n783_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n232_), .B1(new_n826_), .B2(new_n577_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n818_), .A2(new_n622_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n824_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  INV_X1    g629(.A(new_n783_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n577_), .A2(KEYINPUT123), .ZN(new_n833_));
  MUX2_X1   g632(.A(KEYINPUT123), .B(new_n833_), .S(G113gat), .Z(new_n834_));
  OAI211_X1 g633(.A(new_n832_), .B(new_n834_), .C1(new_n825_), .C2(new_n830_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n827_), .A2(new_n835_), .ZN(G1340gat));
  NOR2_X1   g635(.A1(new_n634_), .A2(KEYINPUT60), .ZN(new_n837_));
  MUX2_X1   g636(.A(KEYINPUT60), .B(new_n837_), .S(new_n233_), .Z(new_n838_));
  NAND2_X1  g637(.A1(new_n825_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT124), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n825_), .A2(KEYINPUT124), .A3(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n523_), .B(new_n832_), .C1(new_n825_), .C2(new_n830_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G120gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1341gat));
  OAI21_X1  g645(.A(new_n227_), .B1(new_n826_), .B2(new_n622_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n622_), .A2(new_n227_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n832_), .B(new_n848_), .C1(new_n825_), .C2(new_n830_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1342gat));
  OAI21_X1  g649(.A(new_n228_), .B1(new_n826_), .B2(new_n665_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n605_), .A2(new_n228_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n832_), .B(new_n852_), .C1(new_n825_), .C2(new_n830_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1343gat));
  NAND2_X1  g653(.A1(new_n822_), .A2(new_n824_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n643_), .A2(new_n394_), .A3(new_n658_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n855_), .A2(new_n576_), .A3(new_n252_), .A4(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g657(.A1(new_n855_), .A2(new_n523_), .A3(new_n252_), .A4(new_n856_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g659(.A1(new_n855_), .A2(new_n666_), .A3(new_n252_), .A4(new_n856_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  AND3_X1   g662(.A1(new_n855_), .A2(new_n252_), .A3(new_n856_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n606_), .A2(G162gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT125), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n855_), .A2(new_n252_), .A3(new_n632_), .A4(new_n856_), .ZN(new_n867_));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n864_), .A2(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1347gat));
  NAND3_X1  g668(.A1(new_n643_), .A2(new_n251_), .A3(new_n445_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n829_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G169gat), .B1(new_n872_), .B2(new_n577_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(KEYINPUT62), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(KEYINPUT126), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n829_), .A2(new_n877_), .A3(new_n871_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n576_), .A2(new_n222_), .ZN(new_n880_));
  OAI22_X1  g679(.A1(new_n874_), .A2(new_n875_), .B1(new_n879_), .B2(new_n880_), .ZN(G1348gat));
  NAND3_X1  g680(.A1(new_n876_), .A2(new_n878_), .A3(new_n523_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n870_), .A2(new_n207_), .A3(new_n634_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n882_), .A2(new_n207_), .B1(new_n855_), .B2(new_n883_), .ZN(G1349gat));
  INV_X1    g683(.A(new_n879_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n622_), .A2(new_n217_), .ZN(new_n886_));
  INV_X1    g685(.A(G183gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n829_), .A2(new_n666_), .A3(new_n871_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n885_), .A2(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1350gat));
  NAND3_X1  g688(.A1(new_n876_), .A2(new_n878_), .A3(new_n606_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G190gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n632_), .A2(new_n283_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n879_), .B2(new_n892_), .ZN(G1351gat));
  NOR2_X1   g692(.A1(new_n648_), .A2(new_n423_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n855_), .A2(new_n576_), .A3(new_n252_), .A4(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g695(.A(new_n894_), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n251_), .B(new_n897_), .C1(new_n822_), .C2(new_n824_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT127), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n266_), .A2(new_n267_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n898_), .A2(new_n899_), .A3(new_n523_), .A4(new_n901_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n855_), .A2(new_n523_), .A3(new_n252_), .A4(new_n894_), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT127), .B1(new_n903_), .B2(G204gat), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n900_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n902_), .B1(new_n904_), .B2(new_n905_), .ZN(G1353gat));
  NAND4_X1  g705(.A1(new_n855_), .A2(new_n666_), .A3(new_n252_), .A4(new_n894_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n611_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT63), .B(G211gat), .Z(new_n910_));
  NAND3_X1  g709(.A1(new_n898_), .A2(new_n666_), .A3(new_n910_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1354gat));
  NAND2_X1  g711(.A1(new_n898_), .A2(new_n632_), .ZN(new_n913_));
  INV_X1    g712(.A(G218gat), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n605_), .A2(new_n914_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n913_), .A2(new_n914_), .B1(new_n898_), .B2(new_n915_), .ZN(G1355gat));
endmodule


