//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  XOR2_X1   g002(.A(G85gat), .B(G92gat), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT7), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n206_), .B(new_n207_), .C1(G99gat), .C2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n209_), .B(new_n210_), .C1(KEYINPUT64), .C2(KEYINPUT7), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n208_), .A2(new_n211_), .A3(KEYINPUT66), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT66), .B1(new_n208_), .B2(new_n211_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT6), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n205_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT67), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(new_n211_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n208_), .A2(new_n211_), .A3(KEYINPUT66), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n216_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n204_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT8), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT8), .B1(new_n216_), .B2(new_n220_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n204_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n228_), .B2(new_n204_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n219_), .A2(new_n227_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT10), .B(G99gat), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n210_), .ZN(new_n236_));
  INV_X1    g035(.A(G85gat), .ZN(new_n237_));
  INV_X1    g036(.A(G92gat), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT9), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n234_), .A2(new_n236_), .A3(new_n239_), .A4(new_n216_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n233_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n244_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n241_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(KEYINPUT35), .B(new_n203_), .C1(new_n248_), .C2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n233_), .A2(new_n240_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n244_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .A4(new_n247_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G190gat), .B(G218gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(G134gat), .B(G162gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT36), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT75), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n264_));
  NAND4_X1  g063(.A1(new_n251_), .A2(new_n264_), .A3(new_n256_), .A4(new_n260_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT74), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT37), .B1(new_n263_), .B2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n267_), .A2(KEYINPUT37), .A3(new_n262_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G1gat), .ZN(new_n271_));
  INV_X1    g070(.A(G8gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT14), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT76), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n276_), .B(KEYINPUT14), .C1(new_n271_), .C2(new_n272_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G1gat), .B(G8gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G231gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT77), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n280_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G57gat), .B(G64gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT68), .B(G71gat), .ZN(new_n286_));
  INV_X1    g085(.A(G78gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n286_), .B(G78gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT11), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n285_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n284_), .B1(new_n288_), .B2(KEYINPUT11), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n283_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G183gat), .B(G211gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G127gat), .B(G155gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT17), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(KEYINPUT79), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n301_), .A2(KEYINPUT17), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n296_), .A2(new_n305_), .A3(new_n302_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT79), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n270_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT80), .ZN(new_n312_));
  XOR2_X1   g111(.A(G197gat), .B(G204gat), .Z(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT21), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G197gat), .B(G204gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT21), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n319_), .A2(KEYINPUT92), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n314_), .A2(new_n315_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(KEYINPUT92), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT23), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(G183gat), .A3(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT22), .B(G169gat), .ZN(new_n331_));
  INV_X1    g130(.A(G176gat), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n328_), .A2(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n334_), .B(KEYINPUT94), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT25), .B(G183gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(KEYINPUT24), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(KEYINPUT24), .A3(new_n334_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n325_), .A2(new_n327_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n344_), .B2(new_n327_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n336_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n323_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT20), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n328_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n352_));
  AOI21_X1  g151(.A(G176gat), .B1(new_n352_), .B2(KEYINPUT22), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G169gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n346_), .B2(new_n329_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n349_), .B1(new_n323_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n348_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT19), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G92gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT18), .B(G64gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n351_), .A2(new_n355_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n368_), .A2(new_n321_), .A3(new_n320_), .A4(new_n322_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n323_), .A2(new_n347_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT20), .A4(new_n360_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n360_), .B1(new_n348_), .B2(new_n357_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n366_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G127gat), .B(G134gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n380_), .B(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G155gat), .A2(G162gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G141gat), .A2(G148gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(KEYINPUT90), .A2(KEYINPUT2), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G141gat), .A2(G148gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(KEYINPUT90), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(new_n389_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n384_), .B(new_n385_), .C1(new_n388_), .C2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT89), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n385_), .B2(KEYINPUT1), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n385_), .A2(KEYINPUT1), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n398_), .A2(KEYINPUT89), .A3(G155gat), .A4(G162gat), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n396_), .A2(new_n397_), .A3(new_n384_), .A4(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n386_), .B(KEYINPUT88), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n390_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n394_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n383_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n376_), .B(new_n378_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n394_), .A2(new_n405_), .A3(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT97), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT97), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n404_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(new_n237_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT0), .B(G57gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT4), .B1(new_n383_), .B2(new_n403_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n409_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n413_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n372_), .A2(new_n375_), .A3(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n404_), .A2(new_n406_), .A3(new_n409_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT95), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n417_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n410_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT96), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT33), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT33), .B1(new_n429_), .B2(new_n430_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n423_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT98), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n426_), .A2(new_n428_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n417_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n429_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n358_), .A2(new_n360_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT99), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT20), .A4(new_n361_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n358_), .A2(KEYINPUT99), .A3(new_n360_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n437_), .B(new_n439_), .C1(new_n445_), .C2(new_n438_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT98), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n423_), .B(new_n447_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n434_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G78gat), .B(G106gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT93), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G50gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n403_), .A2(KEYINPUT29), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n454_), .A2(KEYINPUT28), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(KEYINPUT28), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n403_), .A2(KEYINPUT29), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n323_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G228gat), .A2(G233gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT91), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(G22gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n460_), .A2(new_n462_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n453_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n460_), .A2(new_n462_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n465_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(new_n467_), .A3(new_n452_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n449_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT27), .B(new_n375_), .C1(new_n445_), .C2(new_n366_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n437_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT27), .B1(new_n372_), .B2(new_n375_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n477_), .A2(new_n474_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT100), .ZN(new_n482_));
  INV_X1    g281(.A(new_n375_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n367_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n479_), .B1(new_n485_), .B2(KEYINPUT27), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT100), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n478_), .A4(new_n474_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n476_), .A2(new_n482_), .A3(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n383_), .B(KEYINPUT85), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(new_n356_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G71gat), .B(G99gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n491_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G15gat), .B(G43gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT30), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n495_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n486_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(new_n474_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n500_), .A2(new_n437_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n489_), .A2(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G120gat), .B(G148gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(G204gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT5), .B(G176gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT70), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n295_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n226_), .B1(new_n225_), .B2(KEYINPUT8), .ZN(new_n513_));
  AOI211_X1 g312(.A(KEYINPUT67), .B(new_n218_), .C1(new_n224_), .C2(new_n204_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n216_), .A2(new_n220_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n218_), .A3(new_n204_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT65), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n228_), .A2(new_n229_), .A3(new_n204_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n513_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n240_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n512_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n233_), .A2(new_n295_), .A3(new_n240_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(KEYINPUT69), .A3(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(KEYINPUT69), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n522_), .A2(KEYINPUT12), .A3(new_n523_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT12), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n241_), .A2(new_n530_), .A3(new_n512_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n511_), .B1(new_n528_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT71), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n523_), .A2(KEYINPUT12), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n295_), .B1(new_n233_), .B2(new_n240_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n531_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n526_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n509_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n533_), .A2(new_n534_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n534_), .B1(new_n533_), .B2(new_n542_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n505_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n533_), .A2(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT71), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n533_), .A2(new_n542_), .A3(new_n534_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(KEYINPUT13), .A3(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n280_), .B(new_n249_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n280_), .A2(new_n249_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n280_), .B2(new_n246_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555_));
  MUX2_X1   g354(.A(new_n552_), .B(new_n554_), .S(new_n555_), .Z(new_n556_));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n556_), .B(KEYINPUT81), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n559_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n504_), .A2(new_n551_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n312_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT101), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(new_n271_), .A3(new_n437_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT38), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n551_), .A2(new_n566_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n263_), .A2(new_n267_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT102), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n310_), .ZN(new_n577_));
  NOR4_X1   g376(.A1(new_n573_), .A2(new_n576_), .A3(new_n577_), .A4(new_n504_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G1gat), .B1(new_n579_), .B2(new_n478_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n571_), .A2(new_n580_), .ZN(G1324gat));
  AOI21_X1  g380(.A(new_n272_), .B1(new_n578_), .B2(new_n501_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT39), .Z(new_n583_));
  NAND3_X1  g382(.A1(new_n569_), .A2(new_n272_), .A3(new_n501_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT40), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(G1325gat));
  INV_X1    g386(.A(G15gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n500_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n578_), .B2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n312_), .A2(new_n588_), .A3(new_n589_), .A4(new_n567_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT104), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n591_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n593_), .A2(KEYINPUT104), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n592_), .A2(new_n594_), .A3(new_n595_), .A4(new_n596_), .ZN(G1326gat));
  OAI21_X1  g396(.A(G22gat), .B1(new_n579_), .B2(new_n475_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT42), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n475_), .A2(G22gat), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n599_), .B1(new_n568_), .B2(new_n600_), .ZN(G1327gat));
  AND2_X1   g400(.A1(new_n263_), .A2(new_n267_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n577_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT106), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n567_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(G29gat), .B1(new_n605_), .B2(new_n437_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n449_), .A2(new_n475_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n482_), .A2(new_n488_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n500_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n502_), .A2(new_n503_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n270_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT105), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT43), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT105), .B(new_n614_), .C1(new_n504_), .C2(new_n270_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n551_), .A2(new_n310_), .A3(new_n566_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT44), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n619_), .A2(G29gat), .A3(new_n437_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n613_), .A2(KEYINPUT44), .A3(new_n615_), .A4(new_n616_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n606_), .B1(new_n620_), .B2(new_n621_), .ZN(G1328gat));
  INV_X1    g421(.A(G36gat), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n621_), .A2(new_n501_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(new_n619_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n605_), .A2(KEYINPUT45), .A3(new_n623_), .A4(new_n501_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT45), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n567_), .A2(new_n623_), .A3(new_n604_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n628_), .B2(new_n486_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT107), .B1(new_n625_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT46), .ZN(new_n632_));
  INV_X1    g431(.A(new_n619_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n621_), .A2(new_n501_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G36gat), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n630_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n631_), .A2(new_n632_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT108), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n635_), .A2(new_n636_), .A3(KEYINPUT46), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n631_), .A2(new_n638_), .A3(KEYINPUT108), .A4(new_n632_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n641_), .A2(new_n642_), .A3(new_n643_), .ZN(G1329gat));
  NAND4_X1  g443(.A1(new_n619_), .A2(G43gat), .A3(new_n589_), .A4(new_n621_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n605_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n500_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(G43gat), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT47), .ZN(G1330gat));
  AND3_X1   g448(.A1(new_n619_), .A2(new_n474_), .A3(new_n621_), .ZN(new_n650_));
  INV_X1    g449(.A(G50gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n474_), .A2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT109), .Z(new_n653_));
  OAI22_X1  g452(.A1(new_n650_), .A2(new_n651_), .B1(new_n646_), .B2(new_n653_), .ZN(G1331gat));
  NOR2_X1   g453(.A1(new_n576_), .A2(new_n504_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n550_), .A2(new_n565_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n310_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(G57gat), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n478_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n504_), .A2(new_n550_), .A3(new_n565_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n312_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n437_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(KEYINPUT110), .A3(new_n658_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT110), .B1(new_n663_), .B2(new_n658_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n659_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT111), .Z(G1332gat));
  OAI21_X1  g467(.A(G64gat), .B1(new_n657_), .B2(new_n486_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT48), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n486_), .A2(G64gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n661_), .B2(new_n671_), .ZN(G1333gat));
  OR3_X1    g471(.A1(new_n661_), .A2(G71gat), .A3(new_n500_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G71gat), .B1(new_n657_), .B2(new_n500_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT112), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT49), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT49), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1334gat));
  OAI21_X1  g477(.A(G78gat), .B1(new_n657_), .B2(new_n475_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n662_), .A2(new_n287_), .A3(new_n474_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1335gat));
  NAND4_X1  g482(.A1(new_n613_), .A2(new_n577_), .A3(new_n615_), .A4(new_n656_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n478_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n660_), .A2(new_n604_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n237_), .A3(new_n437_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT114), .ZN(G1336gat));
  OAI21_X1  g489(.A(G92gat), .B1(new_n684_), .B2(new_n486_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n687_), .A2(new_n238_), .A3(new_n501_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT115), .ZN(G1337gat));
  OAI21_X1  g493(.A(G99gat), .B1(new_n684_), .B2(new_n500_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n235_), .A3(new_n589_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g497(.A1(new_n687_), .A2(new_n210_), .A3(new_n474_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n684_), .A2(new_n475_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT52), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(G106gat), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n700_), .B2(G106gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n699_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR4_X1   g505(.A1(new_n501_), .A2(new_n500_), .A3(new_n478_), .A4(new_n474_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT55), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n539_), .A2(KEYINPUT117), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT117), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT55), .B1(new_n532_), .B2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n529_), .A2(new_n527_), .A3(new_n531_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n511_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT119), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n511_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT56), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT119), .B(KEYINPUT56), .C1(new_n714_), .C2(new_n511_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n715_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n552_), .A2(new_n555_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n554_), .B(KEYINPUT118), .Z(new_n723_));
  OAI211_X1 g522(.A(new_n559_), .B(new_n722_), .C1(new_n723_), .C2(new_n555_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n562_), .A2(new_n542_), .A3(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n721_), .A2(KEYINPUT58), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT58), .B1(new_n721_), .B2(new_n725_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n270_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n565_), .A2(new_n542_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT56), .B1(new_n714_), .B2(new_n511_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n731_), .B2(new_n715_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n562_), .A2(new_n724_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n574_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT57), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n511_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n542_), .B(new_n565_), .C1(new_n738_), .C2(new_n730_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n734_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(KEYINPUT57), .A3(new_n574_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n737_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n577_), .B1(new_n728_), .B2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n545_), .A2(new_n549_), .A3(new_n310_), .A4(new_n566_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT116), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n746_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n270_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT54), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n550_), .A2(KEYINPUT116), .A3(new_n310_), .A4(new_n566_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n745_), .A2(new_n746_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n270_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n750_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n708_), .B1(new_n744_), .B2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G113gat), .B1(new_n757_), .B2(new_n565_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT120), .Z(new_n759_));
  XOR2_X1   g558(.A(new_n707_), .B(KEYINPUT121), .Z(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(KEYINPUT59), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n754_), .B1(new_n753_), .B2(new_n270_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n268_), .A2(new_n269_), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT54), .B(new_n763_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  AOI211_X1 g564(.A(new_n736_), .B(new_n602_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT57), .B1(new_n741_), .B2(new_n574_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n721_), .A2(new_n725_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n721_), .A2(KEYINPUT58), .A3(new_n725_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n763_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n310_), .B1(new_n768_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n761_), .B1(new_n765_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT59), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n757_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT122), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n775_), .B(KEYINPUT122), .C1(new_n757_), .C2(new_n776_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n565_), .A2(G113gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n759_), .B1(new_n781_), .B2(new_n782_), .ZN(G1340gat));
  OR2_X1    g582(.A1(new_n777_), .A2(new_n550_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT60), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n550_), .B2(G120gat), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n757_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G120gat), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1341gat));
  AOI21_X1  g589(.A(G127gat), .B1(new_n757_), .B2(new_n310_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n310_), .A2(G127gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n781_), .B2(new_n792_), .ZN(G1342gat));
  INV_X1    g592(.A(G134gat), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n270_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n779_), .A2(new_n780_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n757_), .A2(new_n576_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n794_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n796_), .A2(KEYINPUT123), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT123), .B1(new_n796_), .B2(new_n798_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1343gat));
  OAI21_X1  g600(.A(new_n437_), .B1(new_n765_), .B2(new_n774_), .ZN(new_n802_));
  NOR4_X1   g601(.A1(new_n802_), .A2(new_n589_), .A3(new_n475_), .A4(new_n501_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n565_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n551_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n310_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT61), .B(G155gat), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  AOI21_X1  g609(.A(G162gat), .B1(new_n803_), .B2(new_n576_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n763_), .A2(G162gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n803_), .B2(new_n812_), .ZN(G1347gat));
  AOI21_X1  g612(.A(new_n474_), .B1(new_n744_), .B2(new_n756_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n500_), .A2(new_n486_), .A3(new_n437_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(new_n331_), .A3(new_n565_), .A4(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n565_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT124), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n819_), .A2(G169gat), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n819_), .B2(G169gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n816_), .B1(new_n821_), .B2(new_n822_), .ZN(G1348gat));
  NAND2_X1  g622(.A1(new_n814_), .A2(new_n815_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n550_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(new_n332_), .ZN(G1349gat));
  NOR3_X1   g625(.A1(new_n824_), .A2(new_n577_), .A3(new_n337_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n827_), .A2(KEYINPUT126), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(KEYINPUT126), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n824_), .A2(new_n577_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(G183gat), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n828_), .A2(new_n829_), .A3(new_n831_), .ZN(G1350gat));
  OAI21_X1  g631(.A(G190gat), .B1(new_n824_), .B2(new_n270_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n576_), .A2(new_n338_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n824_), .B2(new_n834_), .ZN(G1351gat));
  AOI211_X1 g634(.A(new_n437_), .B(new_n475_), .C1(new_n744_), .C2(new_n756_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n589_), .A2(new_n486_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n565_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n551_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g642(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n310_), .A2(new_n844_), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT127), .Z(new_n846_));
  NOR2_X1   g645(.A1(new_n838_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1354gat));
  AND3_X1   g648(.A1(new_n839_), .A2(G218gat), .A3(new_n763_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G218gat), .B1(new_n839_), .B2(new_n576_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1355gat));
endmodule


