//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n978_, new_n979_, new_n981_, new_n982_, new_n984_, new_n985_,
    new_n986_, new_n988_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_;
  INV_X1    g000(.A(KEYINPUT33), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT86), .ZN(new_n203_));
  INV_X1    g002(.A(G134gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G127gat), .ZN(new_n205_));
  INV_X1    g004(.A(G127gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G134gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n208_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n211_));
  INV_X1    g010(.A(G120gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G113gat), .ZN(new_n213_));
  INV_X1    g012(.A(G113gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G120gat), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT85), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT85), .B1(new_n213_), .B2(new_n215_), .ZN(new_n217_));
  OAI22_X1  g016(.A1(new_n210_), .A2(new_n211_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n206_), .A2(G134gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n204_), .A2(G127gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT84), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT85), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n214_), .A2(G120gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n212_), .A2(G113gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT85), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n221_), .A2(new_n225_), .A3(new_n209_), .A4(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n203_), .B1(new_n218_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G141gat), .ZN(new_n229_));
  INV_X1    g028(.A(G148gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G155gat), .B(G162gat), .Z(new_n235_));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n238_), .A2(KEYINPUT88), .B1(G141gat), .B2(G148gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT88), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT2), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n239_), .A2(new_n241_), .B1(new_n231_), .B2(KEYINPUT3), .ZN(new_n242_));
  NAND3_X1  g041(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT89), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(KEYINPUT89), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT87), .B1(new_n231_), .B2(KEYINPUT3), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n242_), .A2(new_n247_), .A3(new_n248_), .A4(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n237_), .B1(new_n252_), .B2(new_n235_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n210_), .A2(new_n211_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n216_), .A2(new_n217_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT86), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n228_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n218_), .A2(new_n227_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT4), .B1(new_n257_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(KEYINPUT86), .ZN(new_n264_));
  INV_X1    g063(.A(new_n256_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n238_), .A2(KEYINPUT88), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n241_), .A2(new_n266_), .A3(new_n233_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n231_), .A2(KEYINPUT3), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n248_), .A2(new_n267_), .A3(new_n268_), .A4(new_n251_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n247_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n235_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n237_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n264_), .A2(new_n265_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n261_), .A2(new_n263_), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n263_), .B1(new_n274_), .B2(new_n259_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(G85gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G57gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n202_), .B1(new_n280_), .B2(new_n285_), .ZN(new_n286_));
  AOI211_X1 g085(.A(KEYINPUT33), .B(new_n284_), .C1(new_n277_), .C2(new_n279_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n263_), .B1(new_n261_), .B2(new_n276_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n274_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n284_), .ZN(new_n290_));
  OAI22_X1  g089(.A1(new_n286_), .A2(new_n287_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  OAI211_X1 g093(.A(KEYINPUT21), .B(new_n292_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT21), .ZN(new_n296_));
  XOR2_X1   g095(.A(G211gat), .B(G218gat), .Z(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(KEYINPUT91), .ZN(new_n298_));
  XOR2_X1   g097(.A(G197gat), .B(G204gat), .Z(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(KEYINPUT21), .B2(new_n293_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n295_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(KEYINPUT24), .A3(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT25), .B(G183gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT26), .B(G190gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n309_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n306_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT78), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n314_), .B(new_n306_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n304_), .A2(KEYINPUT24), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(KEYINPUT23), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n320_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(KEYINPUT23), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n316_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n313_), .A2(new_n315_), .A3(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n320_), .A2(G183gat), .A3(G190gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(new_n326_), .A3(KEYINPUT81), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n318_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n328_));
  INV_X1    g127(.A(G183gat), .ZN(new_n329_));
  INV_X1    g128(.A(G190gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT82), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT82), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n327_), .A2(new_n328_), .A3(new_n334_), .A4(new_n331_), .ZN(new_n335_));
  AOI21_X1  g134(.A(G176gat), .B1(KEYINPUT80), .B2(KEYINPUT22), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G169gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n302_), .B1(new_n325_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT19), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n323_), .A2(new_n331_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n305_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT22), .B(G169gat), .ZN(new_n345_));
  INV_X1    g144(.A(G176gat), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(KEYINPUT94), .A2(KEYINPUT24), .ZN(new_n349_));
  NOR2_X1   g148(.A1(KEYINPUT94), .A2(KEYINPUT24), .ZN(new_n350_));
  OAI211_X1 g149(.A(KEYINPUT95), .B(new_n305_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n304_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT95), .B1(new_n353_), .B2(new_n305_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n329_), .A2(KEYINPUT25), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G183gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n330_), .A2(KEYINPUT26), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G190gat), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .A4(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n350_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(KEYINPUT94), .A2(KEYINPUT24), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n303_), .A3(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n362_), .A2(new_n365_), .A3(new_n327_), .A4(new_n328_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n348_), .B1(new_n355_), .B2(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT20), .B(new_n342_), .C1(new_n367_), .C2(new_n301_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT96), .B1(new_n339_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n315_), .A2(new_n324_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(KEYINPUT77), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n314_), .B1(new_n373_), .B2(new_n306_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n338_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n301_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT96), .ZN(new_n377_));
  INV_X1    g176(.A(new_n368_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n338_), .B(new_n302_), .C1(new_n370_), .C2(new_n374_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n367_), .B2(new_n301_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n341_), .B(KEYINPUT93), .Z(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT98), .ZN(new_n387_));
  XOR2_X1   g186(.A(KEYINPUT97), .B(KEYINPUT18), .Z(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n369_), .A2(new_n379_), .A3(new_n385_), .A4(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT99), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n368_), .B1(new_n375_), .B2(new_n301_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n395_), .A2(new_n377_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n396_), .A2(KEYINPUT99), .A3(new_n391_), .A4(new_n369_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n369_), .A2(new_n385_), .A3(new_n379_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n391_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT100), .B1(new_n291_), .B2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n288_), .A2(new_n290_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n275_), .B1(new_n274_), .B2(new_n259_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n228_), .A2(new_n256_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT4), .B1(new_n405_), .B2(new_n273_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n404_), .A2(new_n262_), .A3(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n285_), .B1(new_n407_), .B2(new_n278_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT33), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n280_), .A2(new_n202_), .A3(new_n285_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n403_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n394_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT100), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n277_), .A2(new_n284_), .A3(new_n279_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n408_), .A2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n391_), .A2(KEYINPUT32), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n398_), .A2(new_n417_), .ZN(new_n418_));
  AND4_X1   g217(.A1(new_n362_), .A2(new_n365_), .A3(new_n327_), .A4(new_n328_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n305_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT95), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n304_), .A3(new_n351_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n419_), .A2(new_n423_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n381_), .B1(new_n424_), .B2(new_n302_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n342_), .B1(new_n376_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n383_), .A2(new_n384_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT101), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n417_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n429_), .B2(new_n417_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n416_), .B(new_n418_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n402_), .A2(new_n414_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n301_), .B1(new_n253_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G106gat), .ZN(new_n437_));
  INV_X1    g236(.A(G106gat), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n438_), .B(new_n301_), .C1(new_n253_), .C2(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(G78gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n437_), .A2(new_n443_), .A3(new_n439_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(KEYINPUT90), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT28), .B1(new_n273_), .B2(KEYINPUT29), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT28), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n253_), .A2(new_n449_), .A3(new_n435_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G22gat), .B(G50gat), .Z(new_n452_));
  OR2_X1    g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n452_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n447_), .A2(new_n455_), .A3(KEYINPUT92), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n447_), .A2(KEYINPUT92), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT92), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n445_), .A2(new_n458_), .A3(new_n446_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(new_n454_), .A3(new_n453_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n456_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n434_), .A2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n392_), .B(KEYINPUT27), .C1(new_n428_), .C2(new_n391_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n415_), .A3(new_n408_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(new_n461_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n401_), .A2(KEYINPUT102), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT102), .B1(new_n401_), .B2(new_n466_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n465_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT103), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n401_), .A2(new_n466_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT102), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n401_), .A2(KEYINPUT102), .A3(new_n466_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT103), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n465_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n462_), .A2(new_n470_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G227gat), .A2(G233gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G15gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n375_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n481_), .A2(new_n482_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n405_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487_));
  INV_X1    g286(.A(G43gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT31), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n481_), .A2(new_n482_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n405_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n483_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n486_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n490_), .B1(new_n486_), .B2(new_n493_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT104), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n461_), .B(new_n463_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n495_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n486_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n416_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n498_), .B1(new_n499_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n463_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n494_), .A2(new_n495_), .A3(new_n416_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n506_), .A2(KEYINPUT104), .A3(new_n507_), .A4(new_n461_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n478_), .A2(new_n497_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G232gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT34), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT35), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT69), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT65), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G85gat), .B(G92gat), .ZN(new_n522_));
  OR2_X1    g321(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT10), .B(G99gat), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n438_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n525_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n521_), .A2(new_n526_), .A3(new_n528_), .A4(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n522_), .A2(KEYINPUT8), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G99gat), .ZN(new_n534_));
  AND2_X1   g333(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n535_));
  NOR2_X1   g334(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n534_), .B(new_n438_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n537_));
  OAI22_X1  g336(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n533_), .B1(new_n521_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT8), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n519_), .A3(new_n538_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n522_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n531_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G29gat), .B(G36gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G43gat), .B(G50gat), .Z(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G43gat), .B(G50gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n546_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(KEYINPUT15), .A3(new_n551_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n545_), .A2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT70), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT70), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n511_), .A2(KEYINPUT35), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n552_), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n545_), .A2(KEYINPUT71), .A3(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT71), .B1(new_n545_), .B2(new_n562_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n514_), .B1(new_n561_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n567_), .A2(new_n513_), .A3(new_n557_), .A4(new_n560_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT72), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n566_), .A2(new_n574_), .A3(new_n573_), .A4(new_n568_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(KEYINPUT73), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT37), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n577_), .A2(KEYINPUT73), .A3(KEYINPUT37), .A4(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT11), .ZN(new_n586_));
  XOR2_X1   g385(.A(G71gat), .B(G78gat), .Z(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n586_), .A2(new_n587_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n585_), .A2(KEYINPUT11), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n588_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(G1gat), .ZN(new_n593_));
  INV_X1    g392(.A(G8gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT14), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT74), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n597_), .B(KEYINPUT14), .C1(new_n593_), .C2(new_n594_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G15gat), .B(G22gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G1gat), .B(G8gat), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n596_), .A2(new_n601_), .A3(new_n598_), .A4(new_n599_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n592_), .B(new_n605_), .Z(new_n606_));
  AND2_X1   g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT16), .ZN(new_n611_));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT67), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(KEYINPUT17), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n609_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n616_), .B1(KEYINPUT17), .B2(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n584_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n603_), .A2(new_n552_), .A3(new_n604_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n605_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT75), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT75), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n605_), .A2(new_n554_), .A3(new_n627_), .A4(new_n555_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n624_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n605_), .A2(new_n562_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n622_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n623_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT76), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G169gat), .B(G197gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n630_), .A2(new_n634_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n634_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(new_n629_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT5), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n645_), .B(new_n646_), .Z(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT12), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n649_), .B(new_n531_), .C1(new_n540_), .C2(new_n544_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n521_), .A2(new_n539_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n532_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n544_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n530_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n652_), .A2(new_n653_), .B1(new_n521_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n615_), .A2(KEYINPUT12), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n592_), .B(new_n650_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n592_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n545_), .A2(new_n615_), .A3(KEYINPUT12), .A4(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n655_), .A2(new_n592_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n661_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n545_), .A2(new_n658_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n648_), .B1(new_n662_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n662_), .A2(new_n667_), .A3(new_n648_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(KEYINPUT13), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT13), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n664_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n673_), .A2(new_n666_), .A3(new_n647_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n668_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT68), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NOR4_X1   g477(.A1(new_n509_), .A2(new_n621_), .A3(new_n643_), .A4(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(new_n593_), .A3(new_n416_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT105), .Z(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT38), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT38), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n509_), .A2(new_n643_), .A3(new_n676_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n577_), .A2(new_n578_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n620_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G1gat), .B1(new_n688_), .B2(new_n502_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n682_), .A2(new_n683_), .A3(new_n689_), .ZN(G1324gat));
  INV_X1    g489(.A(new_n506_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n679_), .A2(new_n594_), .A3(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n684_), .A2(new_n691_), .A3(new_n687_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G8gat), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT39), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(KEYINPUT39), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n697_), .B(new_n699_), .ZN(G1325gat));
  OAI21_X1  g499(.A(G15gat), .B1(new_n688_), .B2(new_n497_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT41), .Z(new_n702_));
  INV_X1    g501(.A(G15gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n679_), .A2(new_n703_), .A3(new_n496_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1326gat));
  OAI21_X1  g504(.A(G22gat), .B1(new_n688_), .B2(new_n461_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT42), .ZN(new_n707_));
  INV_X1    g506(.A(G22gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n461_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n679_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1327gat));
  NAND2_X1  g510(.A1(new_n478_), .A2(new_n497_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n504_), .A2(new_n508_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n676_), .A2(new_n643_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n577_), .A2(new_n578_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n620_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n714_), .A2(new_n715_), .A3(new_n717_), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n718_), .A2(G29gat), .A3(new_n502_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n509_), .B2(new_n584_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n721_));
  AOI22_X1  g520(.A1(new_n461_), .A2(new_n434_), .B1(new_n469_), .B2(KEYINPUT103), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n496_), .B1(new_n722_), .B2(new_n477_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n504_), .A2(new_n508_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n721_), .B(new_n583_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n720_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n715_), .A2(new_n686_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n730_), .B(new_n727_), .C1(new_n720_), .C2(new_n725_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n416_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G29gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n732_), .B2(new_n416_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n719_), .B1(new_n735_), .B2(new_n736_), .ZN(G1328gat));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n729_), .A2(new_n731_), .A3(new_n506_), .ZN(new_n739_));
  INV_X1    g538(.A(G36gat), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n714_), .A2(new_n715_), .A3(new_n717_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n506_), .A2(G36gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT109), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747_));
  INV_X1    g546(.A(new_n745_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n718_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n743_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n744_), .A2(KEYINPUT109), .A3(new_n745_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n718_), .B2(new_n748_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n742_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n750_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n738_), .B1(new_n741_), .B2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n750_), .A2(new_n753_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(KEYINPUT46), .C1(new_n739_), .C2(new_n740_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1329gat));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n721_), .B1(new_n714_), .B2(new_n583_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n509_), .A2(KEYINPUT43), .A3(new_n584_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n728_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n730_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n726_), .A2(KEYINPUT44), .A3(new_n728_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n497_), .A2(new_n488_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .A4(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n766_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n729_), .A2(new_n731_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n744_), .A2(new_n496_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n764_), .B1(new_n770_), .B2(new_n488_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n759_), .B(new_n767_), .C1(new_n769_), .C2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n763_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n771_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n759_), .B1(new_n776_), .B2(new_n767_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n774_), .A2(new_n777_), .ZN(G1330gat));
  OR3_X1    g577(.A1(new_n718_), .A2(G50gat), .A3(new_n461_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n732_), .A2(KEYINPUT111), .A3(new_n709_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G50gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT111), .B1(new_n732_), .B2(new_n709_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n781_), .B2(new_n782_), .ZN(G1331gat));
  NAND2_X1  g582(.A1(new_n639_), .A2(new_n642_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n509_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n676_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n621_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(G57gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n416_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n620_), .A2(new_n643_), .ZN(new_n792_));
  NOR4_X1   g591(.A1(new_n509_), .A2(new_n685_), .A3(new_n677_), .A4(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n416_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n790_), .B2(new_n794_), .ZN(G1332gat));
  INV_X1    g594(.A(G64gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(new_n793_), .B2(new_n691_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT48), .Z(new_n798_));
  NAND3_X1  g597(.A1(new_n789_), .A2(new_n796_), .A3(new_n691_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1333gat));
  INV_X1    g599(.A(G71gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n793_), .B2(new_n496_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT49), .Z(new_n803_));
  NAND3_X1  g602(.A1(new_n789_), .A2(new_n801_), .A3(new_n496_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1334gat));
  AOI21_X1  g604(.A(new_n442_), .B1(new_n793_), .B2(new_n709_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT50), .Z(new_n807_));
  NAND2_X1  g606(.A1(new_n709_), .A2(new_n442_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n788_), .B2(new_n808_), .ZN(G1335gat));
  INV_X1    g608(.A(G85gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n676_), .A2(new_n686_), .A3(new_n643_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n720_), .B2(new_n725_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n810_), .B1(new_n812_), .B2(new_n416_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n785_), .A2(new_n678_), .A3(new_n717_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n814_), .A2(G85gat), .A3(new_n502_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n813_), .A2(new_n815_), .ZN(G1336gat));
  NOR3_X1   g615(.A1(new_n814_), .A2(G92gat), .A3(new_n506_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n691_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(G92gat), .B2(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT112), .ZN(G1337gat));
  AOI21_X1  g619(.A(new_n534_), .B1(new_n812_), .B2(new_n496_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n814_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n496_), .A2(new_n527_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g624(.A1(new_n822_), .A2(new_n438_), .A3(new_n709_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n812_), .A2(new_n709_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(G106gat), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n438_), .B(new_n827_), .C1(new_n812_), .C2(new_n709_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n826_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT53), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n826_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1339gat));
  INV_X1    g635(.A(new_n792_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n584_), .A2(new_n786_), .A3(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n838_), .B(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n674_), .B2(new_n643_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n670_), .A2(KEYINPUT115), .A3(new_n784_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n657_), .A2(new_n664_), .A3(new_n659_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n662_), .A2(KEYINPUT55), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n673_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n848_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n846_), .B1(new_n852_), .B2(new_n648_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n854_));
  AOI211_X1 g653(.A(KEYINPUT55), .B(new_n664_), .C1(new_n657_), .C2(new_n659_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n847_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(KEYINPUT56), .A3(new_n647_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n845_), .B1(new_n853_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n626_), .A2(new_n628_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(new_n622_), .A3(new_n633_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n638_), .B1(new_n632_), .B2(new_n623_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n639_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n716_), .B1(new_n858_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n843_), .A2(new_n844_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n857_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT56), .B1(new_n856_), .B2(new_n647_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n864_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(KEYINPUT57), .A3(new_n716_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n857_), .A2(KEYINPUT116), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n856_), .A2(new_n876_), .A3(KEYINPUT56), .A4(new_n647_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n877_), .A3(new_n853_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n674_), .A2(new_n863_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(KEYINPUT58), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n583_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT58), .B1(new_n878_), .B2(new_n879_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n867_), .B(new_n874_), .C1(new_n881_), .C2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n686_), .B1(new_n883_), .B2(KEYINPUT117), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n873_), .B2(new_n716_), .ZN(new_n886_));
  AOI211_X1 g685(.A(new_n866_), .B(new_n685_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n878_), .A2(new_n879_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n583_), .A3(new_n880_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n885_), .B1(new_n888_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n841_), .B1(new_n884_), .B2(new_n893_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n499_), .A2(new_n497_), .A3(new_n502_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT118), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT59), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n838_), .A2(new_n840_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n838_), .A2(new_n840_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n899_), .A2(new_n900_), .B1(new_n686_), .B2(new_n883_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n896_), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n901_), .A2(KEYINPUT59), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n898_), .A2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G113gat), .B1(new_n904_), .B2(new_n643_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n883_), .A2(KEYINPUT117), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n892_), .A2(new_n885_), .A3(new_n867_), .A4(new_n874_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(new_n686_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n902_), .B1(new_n908_), .B2(new_n841_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n214_), .A3(new_n784_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n910_), .ZN(G1340gat));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n903_), .B(new_n678_), .C1(new_n909_), .C2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n898_), .A2(KEYINPUT119), .A3(new_n678_), .A4(new_n903_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n916_), .A3(G120gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n212_), .B1(new_n786_), .B2(KEYINPUT60), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n909_), .B(new_n918_), .C1(KEYINPUT60), .C2(new_n212_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1341gat));
  OAI21_X1  g719(.A(G127gat), .B1(new_n904_), .B2(new_n686_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n909_), .A2(new_n206_), .A3(new_n620_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1342gat));
  OAI21_X1  g722(.A(new_n204_), .B1(new_n897_), .B2(new_n716_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(KEYINPUT120), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n904_), .A2(new_n204_), .A3(new_n584_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1343gat));
  NOR2_X1   g726(.A1(new_n496_), .A2(new_n461_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n928_), .A2(new_n416_), .A3(new_n506_), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n894_), .A2(KEYINPUT121), .A3(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(KEYINPUT121), .B1(new_n894_), .B2(new_n929_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n933_), .A2(new_n229_), .A3(new_n784_), .ZN(new_n934_));
  OAI21_X1  g733(.A(G141gat), .B1(new_n932_), .B2(new_n643_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1344gat));
  NAND3_X1  g735(.A1(new_n933_), .A2(new_n230_), .A3(new_n678_), .ZN(new_n937_));
  OAI21_X1  g736(.A(G148gat), .B1(new_n932_), .B2(new_n677_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1345gat));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  OR3_X1    g739(.A1(new_n932_), .A2(new_n686_), .A3(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n932_), .B2(new_n686_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1346gat));
  NAND2_X1  g742(.A1(new_n583_), .A2(G162gat), .ZN(new_n944_));
  XOR2_X1   g743(.A(new_n944_), .B(KEYINPUT123), .Z(new_n945_));
  NOR2_X1   g744(.A1(new_n932_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n894_), .A2(new_n929_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n894_), .A2(KEYINPUT121), .A3(new_n929_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n716_), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  OAI21_X1  g750(.A(KEYINPUT122), .B1(new_n951_), .B2(G162gat), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953_));
  INV_X1    g752(.A(G162gat), .ZN(new_n954_));
  OAI211_X1 g753(.A(new_n953_), .B(new_n954_), .C1(new_n932_), .C2(new_n716_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n946_), .B1(new_n952_), .B2(new_n955_), .ZN(G1347gat));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n691_), .A2(new_n461_), .A3(new_n507_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n901_), .A2(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(new_n784_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n961_));
  AND4_X1   g760(.A1(new_n957_), .A2(new_n960_), .A3(new_n961_), .A4(G169gat), .ZN(new_n962_));
  INV_X1    g761(.A(G169gat), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n963_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n960_), .A2(new_n964_), .B1(new_n957_), .B2(new_n961_), .ZN(new_n965_));
  INV_X1    g764(.A(new_n959_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n784_), .A2(new_n345_), .ZN(new_n967_));
  XOR2_X1   g766(.A(new_n967_), .B(KEYINPUT125), .Z(new_n968_));
  OAI22_X1  g767(.A1(new_n962_), .A2(new_n965_), .B1(new_n966_), .B2(new_n968_), .ZN(G1348gat));
  INV_X1    g768(.A(new_n894_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n970_), .A2(new_n958_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n971_), .A2(G176gat), .A3(new_n678_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973_));
  AND2_X1   g772(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n972_), .A2(new_n973_), .ZN(new_n975_));
  AOI21_X1  g774(.A(G176gat), .B1(new_n959_), .B2(new_n676_), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n974_), .A2(new_n975_), .A3(new_n976_), .ZN(G1349gat));
  AOI21_X1  g776(.A(G183gat), .B1(new_n971_), .B2(new_n620_), .ZN(new_n978_));
  NOR3_X1   g777(.A1(new_n966_), .A2(new_n307_), .A3(new_n686_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n978_), .A2(new_n979_), .ZN(G1350gat));
  OAI21_X1  g779(.A(G190gat), .B1(new_n966_), .B2(new_n584_), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n959_), .A2(new_n308_), .A3(new_n685_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(G1351gat));
  NAND3_X1  g782(.A1(new_n691_), .A2(new_n928_), .A3(new_n502_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n970_), .A2(new_n984_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n985_), .A2(new_n784_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n986_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g786(.A1(new_n985_), .A2(new_n678_), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g788(.A1(new_n985_), .A2(new_n620_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n991_));
  AND2_X1   g790(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n992_));
  NOR3_X1   g791(.A1(new_n990_), .A2(new_n991_), .A3(new_n992_), .ZN(new_n993_));
  AOI21_X1  g792(.A(new_n993_), .B1(new_n990_), .B2(new_n991_), .ZN(G1354gat));
  INV_X1    g793(.A(G218gat), .ZN(new_n995_));
  AOI21_X1  g794(.A(new_n995_), .B1(new_n985_), .B2(new_n583_), .ZN(new_n996_));
  INV_X1    g795(.A(new_n996_), .ZN(new_n997_));
  NOR2_X1   g796(.A1(new_n716_), .A2(G218gat), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n985_), .A2(new_n998_), .ZN(new_n999_));
  NAND3_X1  g798(.A1(new_n997_), .A2(KEYINPUT127), .A3(new_n999_), .ZN(new_n1000_));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n1001_));
  INV_X1    g800(.A(new_n999_), .ZN(new_n1002_));
  OAI21_X1  g801(.A(new_n1001_), .B1(new_n1002_), .B2(new_n996_), .ZN(new_n1003_));
  NAND2_X1  g802(.A1(new_n1000_), .A2(new_n1003_), .ZN(G1355gat));
endmodule


