//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT24), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT76), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT76), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT24), .A4(new_n202_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n205_), .A2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT26), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT75), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n214_), .B(new_n217_), .C1(new_n218_), .C2(KEYINPUT75), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n211_), .A2(new_n219_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G183gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n215_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n230_), .A3(new_n220_), .ZN(new_n231_));
  AND2_X1   g030(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n207_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n234_), .A3(new_n202_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n225_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT30), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G127gat), .B(G134gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G120gat), .ZN(new_n240_));
  INV_X1    g039(.A(G113gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT77), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT77), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G113gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n240_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n244_), .A3(new_n240_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n239_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n247_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n249_), .A2(new_n245_), .A3(new_n238_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n237_), .B(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G15gat), .B(G43gat), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT31), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G71gat), .B(G99gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n254_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n255_), .B2(new_n259_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT93), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(KEYINPUT78), .A2(G141gat), .A3(G148gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G141gat), .ZN(new_n271_));
  INV_X1    g070(.A(G148gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT1), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT79), .ZN(new_n276_));
  INV_X1    g075(.A(G155gat), .ZN(new_n277_));
  INV_X1    g076(.A(G162gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n270_), .B(new_n273_), .C1(new_n275_), .C2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n280_), .A3(new_n274_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT81), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT81), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n279_), .A2(new_n285_), .A3(new_n280_), .A4(new_n274_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n288_), .A2(new_n271_), .A3(new_n272_), .A4(KEYINPUT80), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT80), .ZN(new_n290_));
  OAI22_X1  g089(.A1(new_n290_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293_));
  INV_X1    g092(.A(new_n268_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT78), .B1(G141gat), .B2(G148gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n265_), .A2(KEYINPUT2), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n292_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n282_), .B1(new_n287_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n251_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n297_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(new_n269_), .B2(new_n293_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n284_), .B(new_n286_), .C1(new_n302_), .C2(new_n292_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n303_), .B(new_n282_), .C1(new_n250_), .C2(new_n248_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n304_), .A3(KEYINPUT4), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT90), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT4), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n251_), .A2(new_n299_), .A3(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n305_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n300_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G85gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n311_), .A2(new_n312_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n264_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n311_), .A2(new_n312_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n317_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n311_), .A2(new_n312_), .A3(new_n317_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(KEYINPUT93), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT27), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT18), .B(G64gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(G92gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT86), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n235_), .A2(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n231_), .A2(new_n234_), .A3(KEYINPUT85), .A4(new_n202_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n214_), .A2(new_n218_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n228_), .B(new_n220_), .C1(new_n208_), .C2(KEYINPUT24), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n203_), .A2(new_n204_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n335_), .A2(new_n336_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G204gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G197gat), .ZN(new_n343_));
  INV_X1    g142(.A(G197gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G204gat), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT82), .B1(new_n344_), .B2(G204gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT21), .ZN(new_n348_));
  AND2_X1   g147(.A1(G211gat), .A2(G218gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G211gat), .A2(G218gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n346_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G211gat), .B(G218gat), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n353_), .A2(KEYINPUT21), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n343_), .A2(new_n345_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n355_), .A2(new_n353_), .A3(KEYINPUT21), .A4(new_n347_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n333_), .B1(new_n341_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n231_), .A2(new_n202_), .A3(new_n234_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n361_));
  INV_X1    g160(.A(new_n216_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n215_), .A2(KEYINPUT26), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n212_), .A2(new_n213_), .B1(new_n216_), .B2(KEYINPUT75), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n364_), .A2(new_n365_), .B1(new_n205_), .B2(new_n210_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n360_), .B1(new_n366_), .B2(new_n224_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n359_), .B1(new_n367_), .B2(new_n357_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n224_), .B(new_n337_), .C1(new_n204_), .C2(new_n203_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n202_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT22), .B(G169gat), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n370_), .B1(new_n371_), .B2(new_n207_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT85), .B1(new_n372_), .B2(new_n231_), .ZN(new_n373_));
  AND4_X1   g172(.A1(KEYINPUT85), .A2(new_n231_), .A3(new_n202_), .A4(new_n234_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n369_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n357_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(KEYINPUT86), .A3(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n358_), .A2(new_n368_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n379_), .B(KEYINPUT19), .Z(new_n380_));
  XOR2_X1   g179(.A(new_n380_), .B(KEYINPUT84), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT87), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT87), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n378_), .A2(new_n385_), .A3(new_n382_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n357_), .A2(new_n369_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n335_), .A2(new_n336_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT89), .A3(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n390_), .A2(KEYINPUT20), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT88), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n367_), .B2(new_n357_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n236_), .A2(KEYINPUT88), .A3(new_n376_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n388_), .A2(new_n389_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n391_), .A2(new_n380_), .A3(new_n395_), .A4(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n332_), .B1(new_n387_), .B2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n378_), .A2(new_n385_), .A3(new_n382_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n385_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n332_), .B(new_n399_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n327_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT94), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n387_), .A2(KEYINPUT94), .A3(new_n332_), .A4(new_n399_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n358_), .A2(new_n368_), .A3(new_n377_), .A4(new_n381_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n357_), .A2(new_n369_), .A3(new_n235_), .ZN(new_n410_));
  AOI211_X1 g209(.A(new_n359_), .B(new_n410_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n411_), .B2(new_n380_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n327_), .B1(new_n412_), .B2(new_n331_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n407_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n405_), .A2(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n263_), .A2(new_n326_), .A3(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G22gat), .B(G50gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT28), .B1(new_n299_), .B2(KEYINPUT29), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n357_), .B1(new_n299_), .B2(KEYINPUT29), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT28), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n303_), .A2(new_n420_), .A3(new_n421_), .A4(new_n282_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n418_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n419_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n417_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(G228gat), .B(G233gat), .C1(new_n357_), .C2(KEYINPUT83), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G78gat), .B(G106gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  NAND2_X1  g228(.A1(new_n418_), .A2(new_n422_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n419_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n417_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n423_), .A3(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n426_), .A2(new_n429_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n429_), .B1(new_n426_), .B2(new_n434_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n416_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT95), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n399_), .B(new_n440_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT92), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n387_), .A2(KEYINPUT92), .A3(new_n399_), .A4(new_n440_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n440_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n324_), .A2(new_n323_), .B1(new_n412_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n399_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n331_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n324_), .A2(KEYINPUT33), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT33), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n311_), .A2(new_n451_), .A3(new_n312_), .A4(new_n317_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n305_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n300_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n322_), .A3(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n449_), .A2(new_n453_), .A3(new_n403_), .A4(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n447_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n437_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n320_), .B(new_n325_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n405_), .A3(new_n414_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n439_), .B1(new_n463_), .B2(new_n263_), .ZN(new_n464_));
  AOI211_X1 g263(.A(KEYINPUT95), .B(new_n262_), .C1(new_n459_), .C2(new_n462_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n438_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT64), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT64), .ZN(new_n471_));
  INV_X1    g270(.A(new_n469_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(new_n467_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  INV_X1    g274(.A(G92gat), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n475_), .A2(new_n476_), .A3(KEYINPUT9), .ZN(new_n477_));
  XOR2_X1   g276(.A(KEYINPUT10), .B(G99gat), .Z(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G85gat), .B(G92gat), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT9), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n474_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n474_), .A2(new_n480_), .A3(KEYINPUT65), .A4(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT8), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT66), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n491_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n472_), .A2(new_n467_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n497_));
  INV_X1    g296(.A(G99gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n498_), .A3(new_n479_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(KEYINPUT66), .A3(new_n492_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n490_), .B1(new_n501_), .B2(new_n481_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n481_), .A2(new_n490_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n493_), .A2(new_n494_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n474_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n489_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n502_), .A2(new_n505_), .A3(new_n489_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n488_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G57gat), .B(G64gat), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n512_));
  XOR2_X1   g311(.A(G71gat), .B(G78gat), .Z(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n512_), .A2(new_n513_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n509_), .A2(KEYINPUT12), .A3(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n485_), .B(new_n486_), .C1(new_n502_), .C2(new_n505_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT12), .B1(new_n519_), .B2(new_n517_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n517_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G230gat), .A2(G233gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n518_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n519_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(new_n516_), .ZN(new_n526_));
  OAI211_X1 g325(.A(G230gat), .B(G233gat), .C1(new_n526_), .C2(new_n521_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G120gat), .B(G148gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G176gat), .B(G204gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  NAND3_X1  g331(.A1(new_n524_), .A2(new_n527_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT13), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OR3_X1    g337(.A1(new_n534_), .A2(new_n537_), .A3(new_n535_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT69), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT15), .ZN(new_n543_));
  INV_X1    g342(.A(G29gat), .ZN(new_n544_));
  INV_X1    g343(.A(G36gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G29gat), .A2(G36gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(G43gat), .ZN(new_n549_));
  INV_X1    g348(.A(G43gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n546_), .A2(new_n550_), .A3(new_n547_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(G50gat), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(G50gat), .B1(new_n549_), .B2(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n543_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(KEYINPUT15), .A3(new_n552_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT73), .B(G22gat), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(G15gat), .ZN(new_n559_));
  INV_X1    g358(.A(G1gat), .ZN(new_n560_));
  INV_X1    g359(.A(G8gat), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT14), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(G15gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n559_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G1gat), .B(G8gat), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n559_), .A2(new_n565_), .A3(new_n562_), .A4(new_n563_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n555_), .A2(new_n557_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n553_), .A2(new_n554_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n569_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n567_), .A2(new_n568_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n573_), .B1(new_n577_), .B2(new_n571_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT74), .B1(new_n575_), .B2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n206_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(new_n344_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(KEYINPUT74), .B(new_n582_), .C1(new_n575_), .C2(new_n578_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n525_), .A2(new_n570_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT34), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT35), .Z(new_n590_));
  INV_X1    g389(.A(new_n508_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n487_), .B1(new_n591_), .B2(new_n506_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n555_), .A2(new_n557_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n587_), .B(new_n590_), .C1(new_n592_), .C2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT70), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n509_), .A2(new_n593_), .B1(new_n525_), .B2(new_n570_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(KEYINPUT35), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n595_), .B(new_n596_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(KEYINPUT70), .A3(new_n590_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G134gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n278_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT36), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n599_), .A2(KEYINPUT72), .A3(new_n600_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n603_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n601_), .A2(new_n610_), .A3(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n607_), .B(KEYINPUT71), .Z(new_n615_));
  NAND3_X1  g414(.A1(new_n599_), .A2(new_n600_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(KEYINPUT37), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n576_), .B(new_n517_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT17), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT16), .B(G183gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(G211gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(G127gat), .B(G155gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  OR3_X1    g426(.A1(new_n622_), .A2(new_n623_), .A3(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(KEYINPUT17), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n622_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n618_), .A2(new_n631_), .ZN(new_n632_));
  AND4_X1   g431(.A1(new_n466_), .A2(new_n542_), .A3(new_n586_), .A4(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n560_), .A3(new_n326_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT38), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n612_), .B(KEYINPUT96), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n631_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n586_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n540_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n466_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n326_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G1gat), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n635_), .A2(new_n642_), .ZN(G1324gat));
  NAND3_X1  g442(.A1(new_n633_), .A2(new_n561_), .A3(new_n415_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT97), .ZN(new_n645_));
  INV_X1    g444(.A(new_n415_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G8gat), .B1(new_n640_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT39), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(G1325gat));
  INV_X1    g450(.A(G15gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n633_), .A2(new_n652_), .A3(new_n262_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT98), .ZN(new_n654_));
  OAI21_X1  g453(.A(G15gat), .B1(new_n640_), .B2(new_n263_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT41), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1326gat));
  XOR2_X1   g456(.A(new_n437_), .B(KEYINPUT99), .Z(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G22gat), .B1(new_n640_), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n633_), .A2(new_n662_), .A3(new_n658_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n639_), .A2(new_n631_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n614_), .A2(KEYINPUT101), .A3(new_n617_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT37), .B1(new_n609_), .B2(new_n611_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n617_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n668_), .B1(new_n466_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n618_), .A2(new_n668_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n461_), .A2(new_n405_), .A3(new_n414_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n437_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n447_), .B2(new_n457_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n263_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT95), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n463_), .A2(new_n439_), .A3(new_n263_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n676_), .B1(new_n683_), .B2(new_n438_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n667_), .B1(new_n675_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT44), .B(new_n667_), .C1(new_n675_), .C2(new_n684_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(G29gat), .A3(new_n326_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n466_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n691_), .A2(new_n612_), .A3(new_n665_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n544_), .B1(new_n693_), .B2(new_n641_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n415_), .A3(new_n688_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  OR2_X1    g496(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n692_), .A2(new_n545_), .A3(new_n415_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n699_), .A2(new_n700_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n697_), .B(new_n698_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(G1329gat));
  OAI21_X1  g504(.A(new_n550_), .B1(new_n693_), .B2(new_n263_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n687_), .A2(G43gat), .A3(new_n262_), .A4(new_n688_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(new_n708_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT47), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n713_), .B(new_n706_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1330gat));
  AOI21_X1  g514(.A(G50gat), .B1(new_n692_), .B2(new_n658_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n678_), .A2(G50gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n689_), .B2(new_n717_), .ZN(G1331gat));
  NAND2_X1  g517(.A1(new_n632_), .A2(new_n540_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n719_), .A2(KEYINPUT105), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(KEYINPUT105), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n691_), .A2(new_n586_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(new_n641_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(G57gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n637_), .A3(new_n541_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n641_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(G57gat), .B2(new_n727_), .ZN(G1332gat));
  OAI21_X1  g527(.A(G64gat), .B1(new_n726_), .B2(new_n646_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT48), .ZN(new_n730_));
  OR3_X1    g529(.A1(new_n723_), .A2(G64gat), .A3(new_n646_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT106), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n730_), .A2(new_n734_), .A3(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n726_), .B2(new_n263_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT49), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n723_), .A2(G71gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n263_), .B2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n726_), .B2(new_n659_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n723_), .A2(G78gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n659_), .B2(new_n743_), .ZN(G1335gat));
  INV_X1    g543(.A(new_n631_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(new_n586_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n540_), .B(new_n746_), .C1(new_n675_), .C2(new_n684_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n475_), .A3(new_n641_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n611_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n599_), .A2(KEYINPUT72), .A3(new_n600_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT72), .B1(new_n599_), .B2(new_n600_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n749_), .B1(new_n752_), .B2(new_n607_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n466_), .A2(new_n541_), .A3(new_n753_), .A4(new_n746_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT107), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n475_), .B1(new_n755_), .B2(new_n641_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n757_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n748_), .B1(new_n758_), .B2(new_n759_), .ZN(G1336gat));
  INV_X1    g559(.A(new_n755_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G92gat), .B1(new_n761_), .B2(new_n415_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT109), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT109), .ZN(new_n764_));
  INV_X1    g563(.A(new_n747_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n415_), .A2(G92gat), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT110), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n763_), .A2(new_n764_), .B1(new_n765_), .B2(new_n767_), .ZN(G1337gat));
  NAND3_X1  g567(.A1(new_n761_), .A2(new_n262_), .A3(new_n478_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n765_), .A2(new_n262_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G99gat), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n770_), .B(G99gat), .C1(new_n747_), .C2(new_n263_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n769_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT51), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n769_), .B(new_n777_), .C1(new_n772_), .C2(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n761_), .A2(new_n479_), .A3(new_n678_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n765_), .A2(new_n678_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(G106gat), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n781_), .B(G106gat), .C1(new_n747_), .C2(new_n437_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n780_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT53), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n780_), .B(new_n788_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1339gat));
  NOR3_X1   g589(.A1(new_n263_), .A2(new_n641_), .A3(new_n415_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n523_), .B1(new_n518_), .B2(new_n522_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n524_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n518_), .A2(new_n522_), .A3(KEYINPUT55), .A4(new_n523_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n532_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(KEYINPUT56), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n532_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(KEYINPUT113), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n586_), .A2(new_n533_), .A3(KEYINPUT112), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT112), .B1(new_n586_), .B2(new_n533_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n801_), .A2(new_n804_), .A3(new_n807_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n575_), .A2(new_n578_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n582_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n593_), .A2(new_n576_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n571_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n569_), .A2(new_n572_), .A3(KEYINPUT114), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n574_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n577_), .A2(new_n573_), .A3(new_n571_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n810_), .B1(new_n817_), .B2(new_n582_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n536_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n808_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n612_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT117), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n753_), .B1(new_n808_), .B2(new_n819_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n821_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n792_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n824_), .A2(KEYINPUT117), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n671_), .A2(new_n672_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n799_), .A2(KEYINPUT56), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n534_), .B1(new_n803_), .B2(new_n802_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n818_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT58), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n829_), .A2(new_n830_), .A3(new_n818_), .A4(new_n833_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n828_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n838_), .B(new_n753_), .C1(new_n808_), .C2(new_n819_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n827_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n745_), .B1(new_n826_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n540_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n632_), .A2(new_n638_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT54), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n632_), .A2(new_n845_), .A3(new_n638_), .A4(new_n842_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n437_), .B(new_n791_), .C1(new_n841_), .C2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849_), .B2(new_n586_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n848_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n820_), .A2(new_n612_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT115), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n824_), .B2(new_n821_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n856_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n835_), .A2(new_n836_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n618_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n824_), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n631_), .B1(new_n858_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n844_), .A2(new_n846_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n678_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT59), .B1(new_n866_), .B2(new_n791_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n851_), .B1(new_n853_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n848_), .A2(new_n852_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(KEYINPUT59), .A3(new_n791_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(KEYINPUT118), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n638_), .A2(new_n241_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n850_), .B1(new_n872_), .B2(new_n873_), .ZN(G1340gat));
  OR2_X1    g673(.A1(new_n240_), .A2(KEYINPUT60), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n240_), .B1(new_n842_), .B2(KEYINPUT60), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT119), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n849_), .A2(new_n875_), .A3(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n878_), .A2(KEYINPUT120), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(KEYINPUT120), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n542_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n881_));
  OAI22_X1  g680(.A1(new_n879_), .A2(new_n880_), .B1(new_n881_), .B2(new_n240_), .ZN(G1341gat));
  AOI21_X1  g681(.A(G127gat), .B1(new_n849_), .B2(new_n745_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n745_), .A2(G127gat), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n872_), .B2(new_n884_), .ZN(G1342gat));
  AOI21_X1  g684(.A(G134gat), .B1(new_n849_), .B2(new_n636_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n618_), .A2(G134gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n872_), .B2(new_n887_), .ZN(G1343gat));
  NOR2_X1   g687(.A1(new_n415_), .A2(new_n641_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n262_), .A2(new_n437_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n889_), .B(new_n890_), .C1(new_n841_), .C2(new_n847_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n638_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n271_), .ZN(G1344gat));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n542_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n272_), .ZN(G1345gat));
  NOR2_X1   g694(.A1(new_n891_), .A2(new_n631_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT121), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n896_), .B(new_n898_), .ZN(G1346gat));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900_));
  INV_X1    g699(.A(new_n636_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n891_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(G162gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n674_), .A2(G162gat), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n891_), .A2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n900_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  OAI221_X1 g705(.A(KEYINPUT122), .B1(new_n891_), .B2(new_n904_), .C1(new_n902_), .C2(G162gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1347gat));
  AOI21_X1  g707(.A(new_n646_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n263_), .A2(new_n326_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(new_n910_), .A3(new_n659_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G169gat), .B1(new_n911_), .B2(new_n638_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n911_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n371_), .A3(new_n586_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT62), .B(G169gat), .C1(new_n911_), .C2(new_n638_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n916_), .A3(new_n917_), .ZN(G1348gat));
  OAI21_X1  g717(.A(new_n207_), .B1(new_n911_), .B2(new_n842_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(KEYINPUT123), .B(new_n207_), .C1(new_n911_), .C2(new_n842_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n866_), .A2(KEYINPUT124), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n910_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n415_), .B1(new_n866_), .B2(KEYINPUT124), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n924_), .A2(new_n925_), .A3(new_n542_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n921_), .A2(new_n922_), .B1(new_n926_), .B2(G176gat), .ZN(G1349gat));
  NOR3_X1   g726(.A1(new_n911_), .A2(new_n214_), .A3(new_n631_), .ZN(new_n928_));
  OR3_X1    g727(.A1(new_n924_), .A2(new_n925_), .A3(new_n631_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n229_), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n911_), .B2(new_n828_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n636_), .A2(new_n218_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n911_), .B2(new_n932_), .ZN(G1351gat));
  NAND3_X1  g732(.A1(new_n909_), .A2(new_n461_), .A3(new_n263_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n638_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n344_), .ZN(G1352gat));
  NOR2_X1   g735(.A1(new_n934_), .A2(new_n542_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n342_), .A2(KEYINPUT125), .ZN(new_n938_));
  XOR2_X1   g737(.A(new_n937_), .B(new_n938_), .Z(G1353gat));
  AOI21_X1  g738(.A(new_n631_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n940_));
  XOR2_X1   g739(.A(new_n940_), .B(KEYINPUT126), .Z(new_n941_));
  NOR2_X1   g740(.A1(new_n934_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1354gat));
  NOR2_X1   g743(.A1(new_n934_), .A2(new_n901_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(G218gat), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n934_), .A2(new_n828_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(G218gat), .B2(new_n947_), .ZN(G1355gat));
endmodule


