//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT24), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT23), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n204_), .A2(KEYINPUT24), .A3(new_n212_), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n205_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT77), .B1(new_n206_), .B2(KEYINPUT25), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n215_), .B(new_n216_), .C1(new_n217_), .C2(KEYINPUT77), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(KEYINPUT79), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT79), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n221_), .B(KEYINPUT23), .C1(new_n206_), .C2(new_n207_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n222_), .A3(new_n210_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n206_), .A2(new_n207_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT78), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n202_), .A2(KEYINPUT22), .ZN(new_n229_));
  AOI21_X1  g028(.A(G176gat), .B1(new_n229_), .B2(new_n227_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n212_), .B1(new_n228_), .B2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n219_), .B1(new_n225_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT30), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G71gat), .B(G99gat), .ZN(new_n235_));
  INV_X1    g034(.A(G43gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G15gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n234_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n241_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT81), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT81), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G155gat), .A3(G162gat), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n250_), .A2(new_n252_), .A3(KEYINPUT1), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT1), .B1(new_n250_), .B2(new_n252_), .ZN(new_n254_));
  OAI22_X1  g053(.A1(new_n253_), .A2(new_n254_), .B1(G155gat), .B2(G162gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n256_), .B(KEYINPUT2), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(KEYINPUT82), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(KEYINPUT82), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT3), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n255_), .A2(new_n259_), .B1(new_n261_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT84), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(KEYINPUT29), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT29), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT84), .B1(new_n268_), .B2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274_));
  INV_X1    g073(.A(G197gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(G204gat), .ZN(new_n276_));
  INV_X1    g075(.A(G204gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G197gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(KEYINPUT21), .A3(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT86), .B1(new_n277_), .B2(G197gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT85), .B1(new_n275_), .B2(G204gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT86), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(new_n275_), .A3(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(new_n277_), .A3(G197gat), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .A4(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT21), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n274_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(new_n279_), .B2(KEYINPUT21), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n280_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G228gat), .A2(G233gat), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n271_), .A2(new_n273_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(KEYINPUT87), .ZN(new_n296_));
  INV_X1    g095(.A(new_n280_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n279_), .A2(KEYINPUT21), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(new_n274_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n297_), .B1(new_n299_), .B2(new_n288_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT87), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n296_), .A2(new_n302_), .B1(new_n269_), .B2(KEYINPUT29), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n295_), .B1(new_n293_), .B2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(KEYINPUT89), .A3(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G22gat), .B(G50gat), .Z(new_n307_));
  NAND3_X1  g106(.A1(new_n268_), .A2(new_n272_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n307_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n311_));
  OR3_X1    g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(KEYINPUT89), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n295_), .B(new_n315_), .C1(new_n293_), .C2(new_n303_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n306_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n305_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n304_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n313_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n295_), .B(new_n305_), .C1(new_n293_), .C2(new_n303_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .A4(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n304_), .A2(new_n318_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n321_), .B1(new_n325_), .B2(new_n322_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT27), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT20), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT91), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n226_), .A2(new_n203_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n212_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n208_), .A2(new_n210_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n334_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n337_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n212_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n226_), .B2(new_n203_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(KEYINPUT91), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n213_), .B1(KEYINPUT24), .B2(new_n204_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n217_), .B2(new_n216_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n223_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n333_), .B1(new_n347_), .B2(new_n292_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n228_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n340_), .B1(new_n349_), .B2(new_n230_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n223_), .B1(G183gat), .B2(G190gat), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n350_), .A2(new_n351_), .B1(new_n218_), .B2(new_n214_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n300_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n332_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n332_), .B1(new_n347_), .B2(new_n292_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT20), .B1(new_n352_), .B2(new_n300_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n354_), .A2(new_n357_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n338_), .A2(new_n342_), .B1(new_n345_), .B2(new_n223_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT20), .B1(new_n364_), .B2(new_n300_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n233_), .A2(new_n292_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n331_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n333_), .B1(new_n233_), .B2(new_n292_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n368_), .B(new_n332_), .C1(new_n292_), .C2(new_n347_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n363_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n328_), .B1(new_n362_), .B2(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n365_), .A2(new_n331_), .A3(new_n366_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n339_), .A2(new_n341_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n296_), .A2(new_n302_), .A3(new_n346_), .A4(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n332_), .B1(new_n374_), .B2(new_n368_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n361_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n367_), .A2(new_n363_), .A3(new_n369_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(KEYINPUT27), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n371_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n327_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT0), .ZN(new_n383_));
  INV_X1    g182(.A(G57gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(G85gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n269_), .A2(new_n388_), .A3(new_n245_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n268_), .A2(new_n393_), .A3(new_n245_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n268_), .A2(new_n393_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n244_), .B1(new_n268_), .B2(new_n393_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n394_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n392_), .B1(new_n398_), .B2(KEYINPUT4), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n269_), .A2(KEYINPUT92), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n395_), .A3(new_n244_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n391_), .B1(new_n401_), .B2(new_n394_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n387_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(new_n390_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n387_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n388_), .B1(new_n401_), .B2(new_n394_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n404_), .B(new_n405_), .C1(new_n406_), .C2(new_n392_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n248_), .A2(new_n381_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT94), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT32), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n361_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n361_), .A2(KEYINPUT93), .A3(new_n411_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT93), .B1(new_n361_), .B2(new_n411_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n367_), .A2(new_n416_), .A3(new_n369_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT33), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n407_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n361_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n398_), .A2(new_n391_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n387_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n389_), .A2(new_n390_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n398_), .B2(KEYINPUT4), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n422_), .B(new_n377_), .C1(new_n424_), .C2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n421_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n407_), .A2(new_n420_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n419_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n317_), .A2(new_n323_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n326_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n410_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n362_), .A2(new_n370_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n399_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n436_), .A2(KEYINPUT33), .A3(new_n404_), .A4(new_n405_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n424_), .A2(new_n426_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n429_), .A2(new_n435_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n408_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(KEYINPUT94), .A3(new_n327_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n379_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n408_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n434_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n409_), .B1(new_n446_), .B2(new_n248_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G229gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G36gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G29gat), .ZN(new_n451_));
  INV_X1    g250(.A(G29gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G36gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n453_), .A3(KEYINPUT69), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G43gat), .B(G50gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT69), .B1(new_n451_), .B2(new_n453_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G8gat), .ZN(new_n460_));
  INV_X1    g259(.A(G22gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G15gat), .ZN(new_n462_));
  INV_X1    g261(.A(G15gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G22gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT14), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n466_), .B1(G1gat), .B2(G8gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n460_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(G1gat), .A2(G8gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(G1gat), .A2(G8gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G15gat), .B(G22gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G1gat), .A2(G8gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT14), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n468_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT69), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n452_), .A2(G36gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n450_), .A2(G29gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n456_), .B1(new_n480_), .B2(new_n454_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n459_), .A2(new_n476_), .A3(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n457_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n483_), .A2(new_n484_), .B1(new_n468_), .B2(new_n475_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n449_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT73), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT15), .B1(new_n459_), .B2(new_n481_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT15), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n484_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n476_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n482_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n448_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT73), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n494_), .B(new_n449_), .C1(new_n482_), .C2(new_n485_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G113gat), .B(G141gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT74), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G169gat), .B(G197gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n487_), .A2(new_n493_), .A3(new_n495_), .A4(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT75), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n487_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT76), .ZN(new_n504_));
  INV_X1    g303(.A(new_n499_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n502_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n505_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT76), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n500_), .A2(new_n501_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G64gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G57gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n384_), .A2(G64gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(KEYINPUT11), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n515_), .B1(KEYINPUT11), .B2(new_n522_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n521_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT10), .B(G99gat), .Z(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G85gat), .A2(G92gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(KEYINPUT9), .A3(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n530_), .A2(KEYINPUT9), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT6), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n528_), .A2(new_n531_), .A3(new_n532_), .A4(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n533_), .B(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT66), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT7), .ZN(new_n543_));
  INV_X1    g342(.A(G99gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n527_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n539_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n538_), .B1(new_n542_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G85gat), .B(G92gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT65), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT65), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n529_), .A2(new_n551_), .A3(new_n530_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT8), .B1(new_n548_), .B2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n550_), .A2(new_n552_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT8), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n534_), .A2(new_n545_), .A3(new_n539_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  AOI211_X1 g357(.A(new_n525_), .B(new_n536_), .C1(new_n554_), .C2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n536_), .B1(new_n554_), .B2(new_n558_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n525_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT12), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n545_), .A2(new_n546_), .A3(new_n539_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n546_), .B1(new_n545_), .B2(new_n539_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n534_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n556_), .B1(new_n565_), .B2(new_n555_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n538_), .A2(new_n541_), .A3(new_n540_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n550_), .A2(new_n556_), .A3(new_n552_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n535_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n525_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n559_), .B1(new_n562_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT64), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT67), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n559_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n560_), .A2(new_n561_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT67), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n578_), .A2(new_n580_), .B1(new_n525_), .B2(new_n570_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n576_), .B1(new_n581_), .B2(new_n575_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT5), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n584_), .B(new_n585_), .Z(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n576_), .B(new_n588_), .C1(new_n581_), .C2(new_n575_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(KEYINPUT13), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n447_), .A2(new_n514_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n570_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n459_), .A2(new_n481_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n560_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT34), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT68), .B(KEYINPUT35), .Z(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n598_), .A3(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n601_), .A2(new_n602_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n605_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n609_), .B(KEYINPUT36), .Z(new_n613_));
  NAND2_X1  g412(.A1(new_n606_), .A2(new_n611_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT70), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT70), .B1(new_n606_), .B2(new_n611_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n612_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT37), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n613_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(KEYINPUT37), .A3(new_n612_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n476_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(new_n525_), .ZN(new_n626_));
  XOR2_X1   g425(.A(G127gat), .B(G155gat), .Z(new_n627_));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT71), .B(KEYINPUT16), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(KEYINPUT17), .A3(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n631_), .B(KEYINPUT17), .Z(new_n634_));
  OAI21_X1  g433(.A(new_n633_), .B1(new_n634_), .B2(new_n626_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n623_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT72), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n595_), .A2(new_n638_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n639_), .A2(G1gat), .A3(new_n444_), .ZN(new_n640_));
  XOR2_X1   g439(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n595_), .A2(new_n636_), .A3(new_n618_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n444_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1324gat));
  OAI21_X1  g444(.A(G8gat), .B1(new_n643_), .B2(new_n380_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n380_), .A2(G8gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT96), .B1(new_n639_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n595_), .A2(new_n652_), .A3(new_n638_), .A4(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT39), .B(G8gat), .C1(new_n643_), .C2(new_n380_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n648_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT98), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n648_), .A2(new_n654_), .A3(new_n658_), .A4(new_n655_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n657_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n643_), .B2(new_n248_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT41), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT41), .ZN(new_n666_));
  INV_X1    g465(.A(new_n639_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n248_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n463_), .A3(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n666_), .A3(new_n669_), .ZN(G1326gat));
  XNOR2_X1  g469(.A(new_n433_), .B(KEYINPUT99), .ZN(new_n671_));
  OAI21_X1  g470(.A(G22gat), .B1(new_n643_), .B2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n671_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n667_), .A2(new_n461_), .A3(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n675_), .A3(new_n677_), .ZN(G1327gat));
  INV_X1    g477(.A(new_n618_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n635_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n595_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n452_), .B1(new_n682_), .B2(new_n444_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n594_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n514_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n635_), .A3(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT101), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n447_), .B2(new_n623_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n620_), .A2(new_n622_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n441_), .A2(new_n327_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n691_), .A2(new_n410_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n668_), .B1(new_n692_), .B2(new_n442_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n689_), .B(new_n690_), .C1(new_n693_), .C2(new_n409_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n687_), .B1(new_n688_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT44), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(G29gat), .A3(new_n408_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n683_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT103), .Z(G1328gat));
  AOI21_X1  g500(.A(new_n699_), .B1(KEYINPUT44), .B2(new_n695_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n450_), .B1(new_n702_), .B2(new_n379_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n682_), .A2(G36gat), .A3(new_n380_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT45), .ZN(new_n706_));
  OR3_X1    g505(.A1(new_n703_), .A2(new_n704_), .A3(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  OAI21_X1  g508(.A(new_n236_), .B1(new_n682_), .B2(new_n248_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT104), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n702_), .A2(G43gat), .A3(new_n668_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(G1330gat));
  INV_X1    g514(.A(new_n682_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G50gat), .B1(new_n716_), .B2(new_n676_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n696_), .A2(G50gat), .A3(new_n433_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n699_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(G1331gat));
  NOR2_X1   g519(.A1(new_n684_), .A2(new_n685_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n693_), .B2(new_n409_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(new_n638_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n384_), .A3(new_n408_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n722_), .A2(new_n635_), .A3(new_n679_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n408_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n727_), .B2(new_n384_), .ZN(G1332gat));
  AOI21_X1  g527(.A(new_n517_), .B1(new_n726_), .B2(new_n379_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n379_), .A2(new_n517_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT107), .Z(new_n733_));
  NAND2_X1  g532(.A1(new_n724_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(G1333gat));
  INV_X1    g534(.A(G71gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n726_), .B2(new_n668_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT49), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n724_), .A2(new_n736_), .A3(new_n668_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n726_), .B2(new_n676_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT50), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n724_), .A2(new_n741_), .A3(new_n676_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n722_), .A2(new_n680_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n408_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT108), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n721_), .A2(new_n635_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n688_), .B2(new_n694_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n444_), .A2(new_n386_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(G1336gat));
  AOI21_X1  g551(.A(G92gat), .B1(new_n746_), .B2(new_n379_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n379_), .A2(G92gat), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT109), .Z(new_n755_));
  AOI21_X1  g554(.A(new_n753_), .B1(new_n750_), .B2(new_n755_), .ZN(G1337gat));
  AOI211_X1 g555(.A(new_n248_), .B(new_n749_), .C1(new_n688_), .C2(new_n694_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT110), .B1(new_n757_), .B2(new_n544_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n688_), .A2(new_n694_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n749_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n668_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(G99gat), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n746_), .A2(new_n526_), .A3(new_n668_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT111), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767_));
  INV_X1    g566(.A(new_n765_), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n767_), .B(new_n768_), .C1(new_n758_), .C2(new_n763_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT112), .B(KEYINPUT51), .C1(new_n766_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n757_), .A2(KEYINPUT110), .A3(new_n544_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n762_), .B1(new_n761_), .B2(G99gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n765_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n767_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n768_), .B1(new_n758_), .B2(new_n763_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT111), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n771_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n776_), .B2(new_n771_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n770_), .B1(new_n778_), .B2(new_n780_), .ZN(G1338gat));
  NAND2_X1  g580(.A1(new_n750_), .A2(new_n433_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(G106gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT113), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n527_), .B1(new_n750_), .B2(new_n433_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n783_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n785_), .B(new_n788_), .C1(new_n783_), .C2(new_n786_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n746_), .A2(new_n527_), .A3(new_n433_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n514_), .A2(new_n636_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n594_), .B2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n685_), .A2(new_n635_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(KEYINPUT114), .C1(new_n591_), .C2(new_n593_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n623_), .A3(new_n800_), .ZN(new_n801_));
  XOR2_X1   g600(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n802_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n798_), .A2(new_n623_), .A3(new_n800_), .A4(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  INV_X1    g607(.A(new_n500_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n491_), .A2(new_n492_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT118), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n449_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n482_), .A2(new_n485_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n499_), .B1(new_n813_), .B2(new_n448_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n809_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n590_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n508_), .A2(new_n513_), .A3(new_n589_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n508_), .A2(new_n513_), .A3(KEYINPUT116), .A4(new_n589_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n560_), .A2(KEYINPUT12), .A3(new_n561_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n571_), .B1(new_n570_), .B2(new_n525_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n579_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n575_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n573_), .A2(KEYINPUT55), .A3(new_n575_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n827_), .B(new_n559_), .C1(new_n562_), .C2(new_n572_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT117), .B1(new_n831_), .B2(KEYINPUT55), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n576_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n830_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n823_), .B1(new_n836_), .B2(new_n588_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n562_), .A2(new_n572_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n575_), .B1(new_n838_), .B2(new_n579_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(KEYINPUT55), .B2(new_n831_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n833_), .B1(new_n576_), .B2(new_n834_), .ZN(new_n841_));
  AOI211_X1 g640(.A(KEYINPUT117), .B(KEYINPUT55), .C1(new_n573_), .C2(new_n575_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(KEYINPUT56), .A3(new_n586_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n837_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n817_), .B1(new_n822_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n808_), .B1(new_n846_), .B2(new_n679_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n836_), .A2(new_n823_), .A3(new_n588_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT56), .B1(new_n843_), .B2(new_n586_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n820_), .A2(new_n821_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n816_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT57), .A3(new_n618_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n815_), .A2(new_n589_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n845_), .B2(new_n856_), .ZN(new_n857_));
  AOI211_X1 g656(.A(KEYINPUT58), .B(new_n855_), .C1(new_n837_), .C2(new_n844_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n690_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n847_), .A2(new_n853_), .A3(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n807_), .B1(new_n636_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n248_), .A2(new_n381_), .A3(new_n444_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n856_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT58), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n845_), .A2(new_n854_), .A3(new_n856_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n623_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n847_), .B(new_n853_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n869_), .B(new_n690_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n635_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n807_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n874_), .A2(new_n863_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n864_), .B1(new_n875_), .B2(new_n862_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G113gat), .B1(new_n876_), .B2(new_n514_), .ZN(new_n877_));
  INV_X1    g676(.A(G113gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(new_n878_), .A3(new_n685_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1340gat));
  OAI21_X1  g679(.A(G120gat), .B1(new_n876_), .B2(new_n684_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n882_));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n594_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n875_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n886_), .ZN(G1341gat));
  OAI21_X1  g686(.A(G127gat), .B1(new_n876_), .B2(new_n635_), .ZN(new_n888_));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n875_), .A2(new_n889_), .A3(new_n636_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1342gat));
  OAI21_X1  g690(.A(G134gat), .B1(new_n876_), .B2(new_n623_), .ZN(new_n892_));
  INV_X1    g691(.A(G134gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n875_), .A2(new_n893_), .A3(new_n679_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1343gat));
  NAND2_X1  g694(.A1(new_n859_), .A2(KEYINPUT119), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n896_), .A2(new_n871_), .A3(new_n853_), .A4(new_n847_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n806_), .B1(new_n897_), .B2(new_n635_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n248_), .A2(new_n408_), .A3(new_n443_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n685_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n594_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G148gat), .ZN(G1345gat));
  NOR3_X1   g703(.A1(new_n898_), .A2(new_n635_), .A3(new_n899_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT120), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1346gat));
  INV_X1    g707(.A(G162gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n900_), .A2(new_n909_), .A3(new_n679_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n898_), .A2(new_n623_), .A3(new_n899_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n909_), .ZN(new_n912_));
  XOR2_X1   g711(.A(new_n912_), .B(KEYINPUT121), .Z(G1347gat));
  NOR3_X1   g712(.A1(new_n248_), .A2(new_n408_), .A3(new_n380_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n914_), .A2(new_n671_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n861_), .A2(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT123), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(new_n685_), .A3(new_n226_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n916_), .A2(new_n685_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n921_), .A2(new_n922_), .A3(G169gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n921_), .B2(G169gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n920_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n927_), .A2(KEYINPUT62), .A3(new_n923_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n919_), .A2(new_n926_), .A3(new_n928_), .ZN(G1348gat));
  NAND2_X1  g728(.A1(new_n918_), .A2(new_n594_), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n874_), .A2(new_n327_), .A3(new_n914_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n684_), .A2(new_n203_), .ZN(new_n932_));
  AOI22_X1  g731(.A1(new_n930_), .A2(new_n203_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  AOI21_X1  g732(.A(G183gat), .B1(new_n931_), .B2(new_n636_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n635_), .A2(new_n217_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(new_n918_), .B2(new_n935_), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n917_), .B2(new_n623_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n679_), .A2(new_n216_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n917_), .B2(new_n938_), .ZN(G1351gat));
  NOR4_X1   g738(.A1(new_n668_), .A2(new_n408_), .A3(new_n327_), .A4(new_n380_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n941_), .B1(new_n873_), .B2(new_n807_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(new_n514_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(G197gat), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(KEYINPUT124), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n947_), .B1(new_n944_), .B2(G197gat), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n946_), .B1(new_n945_), .B2(new_n948_), .ZN(G1352gat));
  AOI21_X1  g748(.A(KEYINPUT125), .B1(new_n942_), .B2(new_n594_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951_));
  NOR4_X1   g750(.A1(new_n898_), .A2(new_n951_), .A3(new_n684_), .A4(new_n941_), .ZN(new_n952_));
  OAI211_X1 g751(.A(KEYINPUT126), .B(G204gat), .C1(new_n950_), .C2(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n874_), .A2(new_n594_), .A3(new_n940_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n951_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n942_), .A2(KEYINPUT125), .A3(new_n594_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n277_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958_));
  INV_X1    g757(.A(new_n954_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n958_), .B1(new_n959_), .B2(new_n277_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n953_), .B1(new_n957_), .B2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(KEYINPUT127), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963_));
  OAI211_X1 g762(.A(new_n963_), .B(new_n953_), .C1(new_n957_), .C2(new_n960_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(G1353gat));
  NOR2_X1   g764(.A1(new_n943_), .A2(new_n635_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AND2_X1   g766(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n966_), .B1(new_n967_), .B2(new_n968_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n969_), .B1(new_n966_), .B2(new_n967_), .ZN(G1354gat));
  OR3_X1    g769(.A1(new_n943_), .A2(G218gat), .A3(new_n618_), .ZN(new_n971_));
  OAI21_X1  g770(.A(G218gat), .B1(new_n943_), .B2(new_n623_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n971_), .A2(new_n972_), .ZN(G1355gat));
endmodule


