//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_;
  XOR2_X1   g000(.A(G22gat), .B(G50gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT28), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(KEYINPUT1), .B2(new_n209_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n207_), .A2(KEYINPUT2), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n205_), .A2(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(KEYINPUT83), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n218_), .A2(new_n221_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT84), .ZN(new_n226_));
  XOR2_X1   g025(.A(G155gat), .B(G162gat), .Z(new_n227_));
  AND3_X1   g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n214_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT85), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(KEYINPUT85), .B(new_n214_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n204_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  AOI211_X1 g035(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n232_), .C2(new_n233_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n236_), .A2(new_n237_), .A3(KEYINPUT86), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT86), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n216_), .B1(G141gat), .B2(G148gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n207_), .A2(KEYINPUT2), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n224_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n221_), .A2(new_n223_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n227_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT84), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT85), .B1(new_n247_), .B2(new_n214_), .ZN(new_n248_));
  AOI211_X1 g047(.A(new_n231_), .B(new_n213_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n235_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT28), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n234_), .A2(new_n204_), .A3(new_n235_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n239_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n203_), .B1(new_n238_), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT86), .B1(new_n236_), .B2(new_n237_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n239_), .A3(new_n252_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n202_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT21), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT88), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT88), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n260_), .A2(new_n265_), .A3(new_n261_), .A4(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT89), .ZN(new_n268_));
  OR3_X1    g067(.A1(new_n260_), .A2(new_n268_), .A3(new_n261_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G228gat), .A2(G233gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT87), .Z(new_n274_));
  OAI211_X1 g073(.A(new_n272_), .B(new_n274_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n213_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n272_), .B1(new_n235_), .B2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(G228gat), .A3(G233gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G78gat), .B(G106gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n254_), .A2(new_n257_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT90), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n254_), .A2(new_n284_), .A3(KEYINPUT90), .A4(new_n257_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n254_), .A2(new_n257_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n283_), .A2(KEYINPUT91), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT91), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n275_), .A2(new_n278_), .A3(new_n291_), .A4(new_n282_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n290_), .A2(new_n281_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n287_), .A2(new_n288_), .A3(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n267_), .A2(new_n271_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT78), .B(G176gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT22), .B(G169gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT23), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(KEYINPUT23), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT79), .A3(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(KEYINPUT79), .B2(new_n302_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n297_), .B(new_n300_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT26), .B(G190gat), .ZN(new_n308_));
  INV_X1    g107(.A(G183gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT76), .B1(new_n309_), .B2(KEYINPUT25), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT25), .B(G183gat), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n308_), .B(new_n310_), .C1(new_n311_), .C2(KEYINPUT76), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT77), .ZN(new_n313_));
  OR2_X1    g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(KEYINPUT24), .A3(new_n297_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n302_), .A2(new_n303_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n314_), .A2(KEYINPUT24), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n313_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n296_), .A2(new_n307_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n311_), .A2(new_n308_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n315_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT92), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n305_), .A2(new_n318_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n299_), .B(KEYINPUT93), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n298_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n328_), .B(new_n297_), .C1(new_n306_), .C2(new_n317_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n272_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n321_), .A2(new_n331_), .A3(KEYINPUT20), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT19), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n296_), .A2(new_n329_), .A3(new_n326_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n320_), .A2(new_n307_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n272_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n334_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n336_), .A2(new_n338_), .A3(KEYINPUT20), .A4(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n335_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n346_), .A2(KEYINPUT27), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n336_), .A2(KEYINPUT20), .A3(new_n338_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n334_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n321_), .A2(new_n331_), .A3(KEYINPUT20), .A4(new_n339_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n344_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n335_), .A2(new_n340_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n344_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n346_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n357_), .B2(KEYINPUT27), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n295_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G227gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(G15gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G71gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT80), .B(G43gat), .ZN(new_n364_));
  INV_X1    g163(.A(G99gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n363_), .B(new_n366_), .Z(new_n367_));
  XNOR2_X1  g166(.A(new_n337_), .B(KEYINPUT30), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n369_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n367_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n367_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G127gat), .B(G134gat), .Z(new_n375_));
  XOR2_X1   g174(.A(G113gat), .B(G120gat), .Z(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  OR3_X1    g179(.A1(new_n372_), .A2(new_n374_), .A3(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n232_), .A2(new_n233_), .A3(new_n377_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n377_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT94), .B1(new_n276_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n232_), .A2(KEYINPUT94), .A3(new_n233_), .A4(new_n377_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT4), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n384_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n384_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n383_), .A2(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n359_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n390_), .A2(new_n384_), .A3(new_n392_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n388_), .A2(new_n394_), .A3(new_n389_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n401_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n403_), .B2(new_n411_), .ZN(new_n412_));
  NOR4_X1   g211(.A1(new_n393_), .A2(KEYINPUT33), .A3(new_n401_), .A4(new_n395_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n357_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n335_), .A2(new_n340_), .A3(KEYINPUT95), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n345_), .A2(KEYINPUT32), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n415_), .A2(new_n349_), .A3(new_n350_), .A4(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n354_), .A2(KEYINPUT95), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n403_), .A3(new_n402_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n422_), .A2(new_n356_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n295_), .A2(new_n423_), .ZN(new_n424_));
  OAI22_X1  g223(.A1(new_n421_), .A2(new_n295_), .B1(new_n405_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n407_), .B1(new_n425_), .B2(new_n383_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G29gat), .B(G36gat), .Z(new_n427_));
  XOR2_X1   g226(.A(G43gat), .B(G50gat), .Z(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT73), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G15gat), .B(G22gat), .ZN(new_n432_));
  INV_X1    g231(.A(G1gat), .ZN(new_n433_));
  INV_X1    g232(.A(G8gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G1gat), .B(G8gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n431_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G229gat), .A2(G233gat), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n429_), .B(KEYINPUT15), .Z(new_n442_));
  INV_X1    g241(.A(new_n438_), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n431_), .B(new_n443_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(new_n440_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G113gat), .B(G141gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT75), .ZN(new_n449_));
  XOR2_X1   g248(.A(G169gat), .B(G197gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT74), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n447_), .B(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n426_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G57gat), .B(G64gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G71gat), .B(G78gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT11), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(KEYINPUT11), .ZN(new_n459_));
  INV_X1    g258(.A(new_n457_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n456_), .A2(KEYINPUT11), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n458_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT67), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n458_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n464_), .A2(KEYINPUT12), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G85gat), .B(G92gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT64), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(KEYINPUT9), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT10), .B(G99gat), .Z(new_n472_));
  INV_X1    g271(.A(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  INV_X1    g274(.A(G92gat), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT9), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(new_n468_), .B2(KEYINPUT64), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n471_), .A2(new_n474_), .A3(new_n478_), .A4(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n365_), .A3(new_n473_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n468_), .A2(KEYINPUT8), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT65), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(KEYINPUT65), .A3(new_n489_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n486_), .A2(new_n487_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n486_), .A2(KEYINPUT66), .A3(new_n487_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n483_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n495_), .B1(new_n500_), .B2(new_n469_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n484_), .B1(new_n494_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n467_), .A2(new_n502_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n496_), .A2(new_n497_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n468_), .B1(new_n504_), .B2(new_n499_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n492_), .B(new_n493_), .C1(new_n505_), .C2(new_n495_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(new_n463_), .A3(new_n484_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n463_), .B1(new_n506_), .B2(new_n484_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n503_), .B(new_n507_), .C1(KEYINPUT12), .C2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G230gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT68), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n484_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n501_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n493_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT65), .B1(new_n488_), .B2(new_n489_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n513_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n464_), .A2(KEYINPUT12), .A3(new_n466_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n507_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n522_));
  INV_X1    g321(.A(new_n463_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT12), .B1(new_n502_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n521_), .A2(new_n522_), .A3(new_n525_), .A4(new_n510_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n512_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n507_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n511_), .B1(new_n528_), .B2(new_n508_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT5), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n527_), .A2(new_n529_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n534_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n537_));
  AND2_X1   g336(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n538_));
  OR3_X1    g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n540_));
  OAI22_X1  g339(.A1(new_n536_), .A2(new_n537_), .B1(new_n540_), .B2(new_n538_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n438_), .B(new_n463_), .ZN(new_n544_));
  AND2_X1   g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G127gat), .B(G155gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(G183gat), .B(G211gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(KEYINPUT67), .A3(KEYINPUT17), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(KEYINPUT17), .B2(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n546_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n502_), .A2(new_n429_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n442_), .A2(new_n502_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT34), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  OAI22_X1  g367(.A1(new_n568_), .A2(KEYINPUT70), .B1(new_n561_), .B2(new_n564_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(KEYINPUT70), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n572_));
  XOR2_X1   g371(.A(G134gat), .B(G162gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n572_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n575_), .A2(new_n572_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n571_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n577_), .B(new_n578_), .C1(new_n579_), .C2(new_n569_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(KEYINPUT71), .A2(KEYINPUT37), .ZN(new_n582_));
  OR2_X1    g381(.A1(KEYINPUT71), .A2(KEYINPUT37), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n576_), .A2(new_n580_), .A3(KEYINPUT71), .A4(KEYINPUT37), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NOR4_X1   g385(.A1(new_n455_), .A2(new_n543_), .A3(new_n558_), .A4(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n587_), .A2(new_n433_), .A3(new_n405_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT38), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n581_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n426_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n543_), .A2(new_n453_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n557_), .A3(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n404_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n589_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n590_), .A2(new_n595_), .A3(new_n596_), .ZN(G1324gat));
  OAI21_X1  g396(.A(G8gat), .B1(new_n594_), .B2(new_n423_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT39), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n587_), .A2(new_n434_), .A3(new_n358_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT96), .B(KEYINPUT40), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1325gat));
  OAI21_X1  g403(.A(G15gat), .B1(new_n594_), .B2(new_n383_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT41), .Z(new_n606_));
  AND2_X1   g405(.A1(new_n381_), .A2(new_n382_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n587_), .A2(new_n361_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(G1326gat));
  INV_X1    g408(.A(new_n295_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G22gat), .B1(new_n594_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT42), .ZN(new_n612_));
  INV_X1    g411(.A(new_n587_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(G22gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT97), .Z(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n613_), .B2(new_n615_), .ZN(G1327gat));
  AND3_X1   g415(.A1(new_n295_), .A2(new_n404_), .A3(new_n423_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n295_), .B1(new_n420_), .B2(new_n414_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n383_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n359_), .A2(new_n406_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n453_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n581_), .A2(new_n557_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n543_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(new_n622_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n405_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n593_), .A2(new_n558_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n621_), .B2(new_n586_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n584_), .A2(new_n585_), .ZN(new_n633_));
  AOI211_X1 g432(.A(KEYINPUT43), .B(new_n633_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT44), .B(new_n630_), .C1(new_n632_), .C2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT43), .B1(new_n426_), .B2(new_n633_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n621_), .A2(new_n631_), .A3(new_n586_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n640_), .A2(KEYINPUT98), .A3(KEYINPUT44), .A4(new_n630_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n630_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n405_), .A2(G29gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n628_), .B1(new_n646_), .B2(new_n647_), .ZN(G1328gat));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT46), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT101), .Z(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(G36gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n423_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n642_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n423_), .A2(G36gat), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n454_), .A2(new_n656_), .A3(new_n625_), .A4(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n657_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT99), .B1(new_n626_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT45), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n658_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n664_));
  OAI22_X1  g463(.A1(new_n663_), .A2(new_n664_), .B1(new_n649_), .B2(KEYINPUT46), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n652_), .B1(new_n655_), .B2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n649_), .A2(KEYINPUT46), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n658_), .A2(new_n660_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT45), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n669_), .B2(new_n662_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n629_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n358_), .B1(new_n671_), .B2(KEYINPUT44), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n637_), .B2(new_n641_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n670_), .B(new_n651_), .C1(new_n673_), .C2(new_n653_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n666_), .A2(new_n674_), .ZN(G1329gat));
  NAND4_X1  g474(.A1(new_n642_), .A2(new_n645_), .A3(G43gat), .A4(new_n607_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G43gat), .B1(new_n627_), .B2(new_n607_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT47), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT47), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(new_n681_), .A3(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1330gat));
  INV_X1    g482(.A(G50gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n627_), .A2(new_n684_), .A3(new_n295_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n610_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n642_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n688_), .B2(G50gat), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT102), .B(new_n684_), .C1(new_n642_), .C2(new_n687_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n689_), .B2(new_n690_), .ZN(G1331gat));
  NAND4_X1  g490(.A1(new_n592_), .A2(new_n453_), .A3(new_n543_), .A4(new_n557_), .ZN(new_n692_));
  INV_X1    g491(.A(G57gat), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n404_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n426_), .B2(new_n622_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n621_), .A2(KEYINPUT103), .A3(new_n453_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n698_), .A2(new_n543_), .A3(new_n557_), .A4(new_n633_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n404_), .B1(new_n699_), .B2(KEYINPUT104), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n700_), .B1(KEYINPUT104), .B2(new_n699_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n694_), .B1(new_n701_), .B2(new_n693_), .ZN(G1332gat));
  OAI21_X1  g501(.A(G64gat), .B1(new_n692_), .B2(new_n423_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT48), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n423_), .A2(G64gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n699_), .B2(new_n705_), .ZN(G1333gat));
  OAI21_X1  g505(.A(G71gat), .B1(new_n692_), .B2(new_n383_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT49), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n383_), .A2(G71gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n699_), .B2(new_n709_), .ZN(G1334gat));
  OAI21_X1  g509(.A(G78gat), .B1(new_n692_), .B2(new_n610_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n610_), .A2(G78gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n699_), .B2(new_n714_), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n542_), .A2(new_n624_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n698_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n475_), .B1(new_n717_), .B2(new_n404_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n542_), .A2(new_n622_), .A3(new_n557_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n640_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n405_), .A2(G85gat), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT106), .Z(new_n723_));
  OAI21_X1  g522(.A(new_n718_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT107), .Z(G1336gat));
  OAI21_X1  g524(.A(G92gat), .B1(new_n721_), .B2(new_n423_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n358_), .A2(new_n476_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n717_), .B2(new_n727_), .ZN(G1337gat));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n607_), .A2(new_n472_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n717_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n720_), .A2(new_n607_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(G99gat), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(G1338gat));
  NAND4_X1  g534(.A1(new_n698_), .A2(new_n473_), .A3(new_n295_), .A4(new_n716_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n640_), .A2(new_n295_), .A3(new_n719_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(G106gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G106gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g541(.A1(new_n610_), .A2(new_n607_), .A3(new_n405_), .A4(new_n423_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT117), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n743_), .A2(KEYINPUT117), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n520_), .A2(new_n524_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n510_), .A2(KEYINPUT111), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n509_), .B1(new_n751_), .B2(new_n510_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n752_), .B2(new_n749_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n512_), .B2(new_n526_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT110), .B(new_n754_), .C1(new_n512_), .C2(new_n526_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n533_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT58), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT115), .ZN(new_n763_));
  NOR2_X1   g562(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n760_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n533_), .B(new_n765_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n440_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n444_), .A2(new_n439_), .A3(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n446_), .A2(new_n767_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n451_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n447_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n451_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n535_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n761_), .A2(new_n763_), .A3(new_n766_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n586_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n773_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n763_), .B1(new_n777_), .B2(new_n766_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  INV_X1    g579(.A(new_n749_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n509_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n748_), .B1(KEYINPUT55), .B2(new_n511_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n781_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n754_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n522_), .B1(new_n748_), .B2(new_n510_), .ZN(new_n786_));
  NOR4_X1   g585(.A1(new_n520_), .A2(new_n524_), .A3(KEYINPUT68), .A4(new_n511_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n784_), .B1(new_n788_), .B2(KEYINPUT110), .ZN(new_n789_));
  INV_X1    g588(.A(new_n758_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n534_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n780_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n759_), .A2(KEYINPUT112), .A3(KEYINPUT56), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n453_), .A2(new_n536_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n772_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT113), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n772_), .B(new_n799_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n796_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n581_), .B1(KEYINPUT116), .B2(KEYINPUT57), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n779_), .B1(new_n806_), .B2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n804_), .B1(new_n796_), .B2(new_n802_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n809_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n557_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n633_), .A2(new_n542_), .A3(new_n453_), .A4(new_n557_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n747_), .B1(new_n814_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n622_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n622_), .A2(new_n535_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n759_), .A2(KEYINPUT112), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n780_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n801_), .B1(new_n824_), .B2(new_n794_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n810_), .B1(new_n825_), .B2(new_n804_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n761_), .A2(new_n766_), .A3(new_n774_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(KEYINPUT115), .A3(new_n762_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n586_), .A3(new_n775_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(new_n813_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n817_), .B1(new_n830_), .B2(new_n558_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n747_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT59), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n829_), .B1(new_n812_), .B2(new_n809_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n825_), .A2(new_n810_), .A3(new_n804_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n558_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n817_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n746_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(KEYINPUT118), .A3(new_n744_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n839_), .A2(new_n846_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n833_), .A2(new_n834_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n834_), .B1(new_n833_), .B2(new_n847_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n453_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n821_), .B1(new_n850_), .B2(new_n820_), .ZN(G1340gat));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n845_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n818_), .B2(KEYINPUT59), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n854_), .B2(new_n543_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n852_), .B1(new_n542_), .B2(KEYINPUT60), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(KEYINPUT120), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n852_), .B2(KEYINPUT60), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n819_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT121), .B1(new_n855_), .B2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n833_), .A2(new_n543_), .A3(new_n847_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G120gat), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n861_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n863_), .A2(new_n867_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n819_), .B2(new_n557_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n848_), .A2(new_n849_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n557_), .A2(G127gat), .ZN(new_n871_));
  XOR2_X1   g670(.A(new_n871_), .B(KEYINPUT122), .Z(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n870_), .B2(new_n872_), .ZN(G1342gat));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n819_), .A2(new_n874_), .A3(new_n591_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n848_), .A2(new_n849_), .A3(new_n633_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n874_), .ZN(G1343gat));
  NOR3_X1   g676(.A1(new_n424_), .A2(new_n607_), .A3(new_n404_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n839_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n622_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n543_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g683(.A1(new_n879_), .A2(KEYINPUT123), .A3(new_n558_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT123), .B1(new_n879_), .B2(new_n558_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n885_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1346gat));
  OR3_X1    g689(.A1(new_n879_), .A2(G162gat), .A3(new_n581_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G162gat), .B1(new_n879_), .B2(new_n633_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1347gat));
  XNOR2_X1  g692(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895_));
  NOR4_X1   g694(.A1(new_n295_), .A2(new_n383_), .A3(new_n405_), .A4(new_n423_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n839_), .A2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n897_), .B2(new_n453_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G169gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n897_), .A2(new_n895_), .A3(new_n453_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n894_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n900_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n894_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n902_), .A2(G169gat), .A3(new_n898_), .A4(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n897_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(new_n327_), .A3(new_n622_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n901_), .A2(new_n904_), .A3(new_n906_), .ZN(G1348gat));
  NOR2_X1   g706(.A1(new_n897_), .A2(new_n542_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n298_), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n908_), .A2(KEYINPUT126), .A3(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT126), .B1(new_n908_), .B2(new_n909_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n908_), .A2(G176gat), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(G1349gat));
  NOR2_X1   g712(.A1(new_n897_), .A2(new_n558_), .ZN(new_n914_));
  MUX2_X1   g713(.A(G183gat), .B(new_n311_), .S(new_n914_), .Z(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n897_), .B2(new_n633_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n591_), .A2(new_n308_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n897_), .B2(new_n917_), .ZN(G1351gat));
  NOR4_X1   g717(.A1(new_n610_), .A2(new_n607_), .A3(new_n405_), .A4(new_n423_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n839_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n622_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n543_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g723(.A1(new_n920_), .A2(new_n557_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  AND2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n928_), .B1(new_n925_), .B2(new_n926_), .ZN(G1354gat));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n920_), .A2(new_n930_), .A3(new_n591_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n839_), .A2(new_n586_), .A3(new_n919_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n931_), .B(KEYINPUT127), .C1(new_n930_), .C2(new_n932_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1355gat));
endmodule


