//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_;
  XNOR2_X1  g000(.A(G71gat), .B(G78gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G57gat), .B(G64gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G57gat), .B(G64gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT11), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n202_), .A3(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT12), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G85gat), .A3(G92gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G85gat), .B(G92gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT10), .B(G99gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G106gat), .ZN(new_n217_));
  OAI221_X1 g016(.A(new_n214_), .B1(new_n215_), .B2(new_n213_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT65), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  NAND3_X1  g024(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n218_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  INV_X1    g030(.A(G99gat), .ZN(new_n232_));
  INV_X1    g031(.A(G106gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n221_), .A2(new_n227_), .A3(new_n230_), .A4(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n215_), .A2(KEYINPUT8), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n224_), .A2(new_n226_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n230_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n234_), .A2(KEYINPUT66), .A3(new_n230_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n215_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n237_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n229_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(KEYINPUT68), .B(new_n237_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT69), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n230_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n240_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n238_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n242_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n215_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n244_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n235_), .A2(new_n236_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n246_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n229_), .ZN(new_n259_));
  AND4_X1   g058(.A1(KEYINPUT69), .A2(new_n258_), .A3(new_n259_), .A4(new_n248_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n212_), .B1(new_n249_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n210_), .B(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n245_), .A2(new_n259_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n264_), .A2(new_n265_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(new_n211_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n261_), .A2(new_n262_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n266_), .ZN(new_n270_));
  OAI211_X1 g069(.A(G230gat), .B(G233gat), .C1(new_n270_), .C2(new_n267_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G120gat), .B(G148gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G204gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G176gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n274_), .B(new_n275_), .Z(new_n276_));
  OR2_X1    g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n276_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(KEYINPUT70), .B2(KEYINPUT13), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT71), .Z(new_n283_));
  NAND2_X1  g082(.A1(G229gat), .A2(G233gat), .ZN(new_n284_));
  INV_X1    g083(.A(G1gat), .ZN(new_n285_));
  INV_X1    g084(.A(G8gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT14), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n285_), .C2(new_n286_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G8gat), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n293_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G29gat), .B(G36gat), .Z(new_n297_));
  XOR2_X1   g096(.A(G43gat), .B(G50gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n294_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT77), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n301_), .A2(KEYINPUT77), .A3(new_n302_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n284_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n299_), .B(KEYINPUT15), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n296_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n309_), .A2(new_n302_), .A3(new_n284_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G113gat), .B(G141gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(G169gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(G197gat), .Z(new_n314_));
  AND3_X1   g113(.A1(new_n311_), .A2(KEYINPUT78), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT78), .B1(new_n311_), .B2(new_n314_), .ZN(new_n316_));
  OAI22_X1  g115(.A1(new_n315_), .A2(new_n316_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n283_), .A2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(G231gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n296_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT74), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n321_), .A2(new_n210_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n210_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G127gat), .B(G155gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT16), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G183gat), .ZN(new_n326_));
  INV_X1    g125(.A(G211gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT17), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n322_), .A2(new_n323_), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n328_), .B(KEYINPUT17), .ZN(new_n332_));
  INV_X1    g131(.A(new_n264_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(new_n320_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n320_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT75), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n332_), .A2(new_n338_), .A3(new_n334_), .A4(new_n335_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT76), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n331_), .A2(new_n337_), .A3(new_n342_), .A4(new_n339_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G78gat), .B(G106gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT92), .Z(new_n347_));
  INV_X1    g146(.A(G233gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT89), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(G228gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(G228gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n348_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G141gat), .B(G148gat), .Z(new_n354_));
  NAND3_X1  g153(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G155gat), .B(G162gat), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n354_), .B(new_n355_), .C1(KEYINPUT1), .C2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT86), .B(KEYINPUT3), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n358_), .A2(G141gat), .A3(G148gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT87), .ZN(new_n360_));
  INV_X1    g159(.A(G141gat), .ZN(new_n361_));
  INV_X1    g160(.A(G148gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT2), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(KEYINPUT2), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n366_));
  AND4_X1   g165(.A1(new_n360_), .A2(new_n364_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n357_), .B1(new_n367_), .B2(new_n356_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n370_), .A2(KEYINPUT21), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G197gat), .B(G204gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(KEYINPUT21), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n370_), .A2(new_n372_), .A3(KEYINPUT21), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n369_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT91), .B1(new_n368_), .B2(KEYINPUT29), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n353_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n368_), .A2(KEYINPUT29), .ZN(new_n381_));
  INV_X1    g180(.A(new_n353_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n377_), .B(KEYINPUT90), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n347_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n347_), .A3(new_n384_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n380_), .A2(new_n384_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n347_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n393_));
  OR3_X1    g192(.A1(new_n368_), .A2(KEYINPUT29), .A3(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G22gat), .B(G50gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n368_), .B2(KEYINPUT29), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n395_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n398_));
  OAI22_X1  g197(.A1(new_n388_), .A2(new_n392_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n400_));
  AND2_X1   g199(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n401_));
  NOR2_X1   g200(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n402_));
  OAI21_X1  g201(.A(G190gat), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n403_), .B(KEYINPUT82), .Z(new_n404_));
  INV_X1    g203(.A(KEYINPUT25), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT26), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(G190gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n410_));
  INV_X1    g209(.A(G183gat), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n405_), .B1(KEYINPUT79), .B2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n404_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G183gat), .A2(G190gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT83), .ZN(new_n416_));
  MUX2_X1   g215(.A(new_n416_), .B(new_n415_), .S(KEYINPUT23), .Z(new_n417_));
  OR2_X1    g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G169gat), .A2(G176gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT24), .A3(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n418_), .A2(KEYINPUT24), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n414_), .A2(new_n417_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(new_n416_), .B2(KEYINPUT23), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT79), .B(G183gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(G190gat), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n419_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT22), .B(G169gat), .ZN(new_n429_));
  INV_X1    g228(.A(G176gat), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n422_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G227gat), .A3(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n433_), .B(KEYINPUT30), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT31), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT31), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n436_), .A2(new_n442_), .A3(new_n439_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G15gat), .B(G43gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT84), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G71gat), .B(G99gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G127gat), .B(G134gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G113gat), .B(G120gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n448_), .B(new_n449_), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n447_), .B(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n441_), .A2(new_n443_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n400_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n389_), .A2(new_n346_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n397_), .A2(new_n398_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n387_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n441_), .A2(new_n443_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n451_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT85), .A3(new_n452_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n399_), .A2(new_n455_), .A3(new_n458_), .A4(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G1gat), .B(G29gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT0), .ZN(new_n465_));
  INV_X1    g264(.A(G57gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G85gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n368_), .A2(new_n450_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n450_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n357_), .B(new_n473_), .C1(new_n367_), .C2(new_n356_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(KEYINPUT4), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT4), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n368_), .A2(new_n476_), .A3(new_n450_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n471_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n472_), .A2(new_n474_), .B1(G225gat), .B2(G233gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n470_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT33), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n482_), .B(new_n470_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n383_), .A2(new_n433_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G226gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT19), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT26), .B(G190gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT25), .B(G183gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n420_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT94), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n424_), .A2(new_n421_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n417_), .B1(G183gat), .B2(G190gat), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n494_), .A2(new_n495_), .B1(new_n496_), .B2(new_n431_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n377_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n486_), .A2(KEYINPUT20), .A3(new_n489_), .A4(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT95), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  OAI221_X1 g301(.A(KEYINPUT20), .B1(new_n497_), .B2(new_n498_), .C1(new_n383_), .C2(new_n433_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n488_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G64gat), .B(G92gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(G8gat), .B(G36gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n475_), .A2(new_n471_), .A3(new_n477_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n472_), .A2(new_n474_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n512_), .B(new_n469_), .C1(new_n471_), .C2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n510_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n502_), .A2(new_n504_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n511_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT97), .B1(new_n485_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n516_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n515_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT97), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n484_), .A4(new_n514_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n478_), .A2(new_n479_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT100), .B1(new_n525_), .B2(new_n469_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n480_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT100), .ZN(new_n528_));
  NOR4_X1   g327(.A1(new_n478_), .A2(new_n528_), .A3(new_n470_), .A4(new_n479_), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n526_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n503_), .A2(new_n488_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n533_));
  NAND2_X1  g332(.A1(new_n499_), .A2(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(KEYINPUT99), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(KEYINPUT99), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n486_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n532_), .B1(new_n537_), .B2(new_n488_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n515_), .A2(KEYINPUT32), .ZN(new_n539_));
  MUX2_X1   g338(.A(new_n538_), .B(new_n505_), .S(new_n539_), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n531_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n463_), .B1(new_n524_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT27), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n516_), .B(KEYINPUT27), .C1(new_n538_), .C2(new_n515_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n530_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n387_), .A2(new_n386_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n389_), .A2(new_n390_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n457_), .B1(new_n549_), .B2(new_n391_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n458_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n455_), .B(new_n462_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n461_), .A2(new_n452_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n399_), .A2(new_n458_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n546_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n345_), .B1(new_n542_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557_));
  XOR2_X1   g356(.A(G134gat), .B(G162gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT36), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n560_), .A2(new_n561_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n308_), .B1(new_n249_), .B2(new_n260_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT72), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT34), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n568_), .A2(KEYINPUT35), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n245_), .A2(new_n299_), .A3(new_n259_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n568_), .A2(KEYINPUT35), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n570_), .A2(new_n565_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n565_), .A2(new_n571_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(new_n574_), .A3(new_n569_), .ZN(new_n575_));
  AOI211_X1 g374(.A(new_n563_), .B(new_n564_), .C1(new_n573_), .C2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n573_), .A2(new_n561_), .A3(new_n560_), .A4(new_n575_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n557_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n564_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n562_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(KEYINPUT37), .A3(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n318_), .A2(new_n556_), .A3(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n285_), .A3(new_n531_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n586_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n576_), .A2(new_n578_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n345_), .B(new_n590_), .C1(new_n542_), .C2(new_n555_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n318_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G1gat), .B1(new_n593_), .B2(new_n530_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n587_), .A2(new_n588_), .A3(new_n594_), .ZN(G1324gat));
  INV_X1    g394(.A(KEYINPUT40), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n544_), .A2(new_n545_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n592_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(G8gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT39), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n601_), .A3(G8gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT102), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n584_), .A2(new_n286_), .A3(new_n597_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n604_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n596_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n608_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(KEYINPUT40), .A3(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(G1325gat));
  INV_X1    g411(.A(G15gat), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n455_), .A2(new_n462_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n592_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n584_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n550_), .A2(new_n551_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n592_), .B2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT42), .Z(new_n623_));
  NAND3_X1  g422(.A1(new_n584_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1327gat));
  NOR2_X1   g424(.A1(new_n590_), .A2(new_n345_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n626_), .B1(new_n542_), .B2(new_n555_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n318_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(G29gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n531_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n583_), .B1(new_n542_), .B2(new_n555_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n345_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n283_), .A2(new_n317_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT43), .B(new_n583_), .C1(new_n542_), .C2(new_n555_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n633_), .A2(new_n634_), .A3(KEYINPUT44), .A4(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT103), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n530_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n629_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n630_), .B1(new_n643_), .B2(new_n644_), .ZN(G1328gat));
  INV_X1    g444(.A(KEYINPUT46), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT106), .ZN(new_n647_));
  INV_X1    g446(.A(new_n627_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n634_), .A2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n650_));
  INV_X1    g449(.A(new_n597_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(G36gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n649_), .A2(new_n650_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n650_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n628_), .B2(new_n652_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n647_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n651_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n637_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n659_), .B2(G36gat), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n646_), .A2(KEYINPUT106), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n661_), .B(new_n657_), .C1(new_n659_), .C2(G36gat), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1329gat));
  INV_X1    g464(.A(new_n637_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n638_), .A2(new_n639_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(G43gat), .A3(new_n553_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n628_), .A2(new_n614_), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n666_), .A2(new_n668_), .B1(G43gat), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g470(.A1(new_n667_), .A2(G50gat), .A3(new_n621_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n649_), .A2(new_n620_), .ZN(new_n673_));
  OAI22_X1  g472(.A1(new_n666_), .A2(new_n672_), .B1(G50gat), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1331gat));
  NOR2_X1   g475(.A1(new_n283_), .A2(new_n317_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n678_), .A2(new_n556_), .A3(new_n583_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G57gat), .B1(new_n679_), .B2(new_n531_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n678_), .A2(new_n591_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n530_), .A2(new_n466_), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n682_), .A2(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(G1332gat));
  INV_X1    g485(.A(G64gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n684_), .B2(new_n597_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT48), .Z(new_n689_));
  NAND3_X1  g488(.A1(new_n679_), .A2(new_n687_), .A3(new_n597_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1333gat));
  INV_X1    g490(.A(G71gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n684_), .B2(new_n614_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT49), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n679_), .A2(new_n692_), .A3(new_n614_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1334gat));
  INV_X1    g495(.A(G78gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n684_), .B2(new_n621_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT50), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n679_), .A2(new_n697_), .A3(new_n621_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1335gat));
  AND2_X1   g500(.A1(new_n633_), .A2(new_n635_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n677_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n530_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n677_), .A2(new_n648_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n531_), .A2(new_n468_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(G1336gat));
  OAI21_X1  g506(.A(G92gat), .B1(new_n703_), .B2(new_n651_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n651_), .A2(G92gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n705_), .B2(new_n709_), .ZN(G1337gat));
  INV_X1    g509(.A(new_n553_), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n705_), .A2(new_n216_), .A3(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n702_), .A2(new_n614_), .A3(new_n677_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(G99gat), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n714_), .B2(G99gat), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n712_), .B(new_n713_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n716_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n723_), .A2(KEYINPUT111), .A3(new_n712_), .A4(new_n713_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n712_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT51), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n721_), .A2(new_n724_), .A3(new_n726_), .ZN(G1338gat));
  NAND4_X1  g526(.A1(new_n633_), .A2(new_n621_), .A3(new_n635_), .A4(new_n677_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G106gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G106gat), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n620_), .A2(new_n217_), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n730_), .A2(new_n731_), .B1(new_n705_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT112), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  OAI221_X1 g534(.A(new_n735_), .B1(new_n705_), .B2(new_n732_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n734_), .A2(KEYINPUT53), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT53), .B1(new_n734_), .B2(new_n736_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1339gat));
  INV_X1    g538(.A(KEYINPUT117), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n305_), .A2(new_n306_), .B1(G229gat), .B2(G233gat), .ZN(new_n741_));
  INV_X1    g540(.A(new_n314_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n309_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n302_), .A2(G229gat), .A3(G233gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n742_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n315_), .A2(new_n316_), .B1(new_n741_), .B2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n261_), .A2(KEYINPUT55), .A3(new_n268_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n262_), .A2(KEYINPUT115), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n748_), .A2(new_n269_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n750_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n261_), .A2(new_n268_), .A3(KEYINPUT55), .A4(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n276_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT56), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n269_), .A2(new_n748_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n749_), .A2(new_n750_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n753_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n276_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n756_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT116), .B(KEYINPUT56), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n755_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n317_), .A2(new_n278_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n747_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n740_), .B1(new_n768_), .B2(new_n589_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT116), .B1(new_n754_), .B2(KEYINPUT56), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT56), .B1(new_n759_), .B2(new_n760_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n756_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n766_), .B1(new_n774_), .B2(new_n755_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT117), .B(new_n590_), .C1(new_n775_), .C2(new_n747_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n769_), .A2(new_n770_), .A3(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT118), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n769_), .A2(new_n776_), .A3(new_n779_), .A4(new_n770_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n768_), .A2(new_n770_), .A3(new_n589_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n746_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n761_), .A2(new_n762_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n772_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI221_X1 g585(.A(new_n782_), .B1(KEYINPUT119), .B2(KEYINPUT58), .C1(new_n783_), .C2(new_n772_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n583_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n781_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n780_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n344_), .B1(new_n778_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n317_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n345_), .A2(KEYINPUT113), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n344_), .B2(new_n317_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n794_), .A2(new_n282_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n583_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT114), .B1(new_n799_), .B2(KEYINPUT54), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n797_), .A2(new_n801_), .A3(new_n802_), .A4(new_n798_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(KEYINPUT54), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n792_), .A2(new_n805_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n554_), .A2(new_n530_), .A3(new_n597_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT59), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n777_), .A2(new_n788_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n811_), .A2(KEYINPUT120), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n781_), .B1(new_n811_), .B2(KEYINPUT120), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n345_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n805_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n810_), .B(new_n807_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n809_), .A2(new_n816_), .A3(new_n317_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G113gat), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n793_), .A2(G113gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n808_), .B2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(new_n283_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n809_), .A2(new_n816_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(KEYINPUT60), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n283_), .B2(KEYINPUT60), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(KEYINPUT121), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(KEYINPUT121), .B2(new_n825_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n822_), .A2(new_n823_), .B1(new_n808_), .B2(new_n827_), .ZN(G1341gat));
  NAND3_X1  g627(.A1(new_n809_), .A2(new_n816_), .A3(new_n345_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G127gat), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n344_), .A2(G127gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n808_), .B2(new_n831_), .ZN(G1342gat));
  NAND3_X1  g631(.A1(new_n809_), .A2(new_n816_), .A3(new_n583_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G134gat), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n590_), .A2(G134gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n808_), .B2(new_n835_), .ZN(G1343gat));
  AOI21_X1  g635(.A(new_n552_), .B1(new_n792_), .B2(new_n805_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n531_), .A3(new_n651_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n793_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(new_n361_), .ZN(G1344gat));
  NOR2_X1   g639(.A1(new_n838_), .A2(new_n283_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n362_), .ZN(G1345gat));
  NOR2_X1   g641(.A1(new_n838_), .A2(new_n344_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT61), .B(G155gat), .Z(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT122), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n843_), .B(new_n845_), .ZN(G1346gat));
  OAI21_X1  g645(.A(G162gat), .B1(new_n838_), .B2(new_n798_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n590_), .A2(G162gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n838_), .B2(new_n848_), .ZN(G1347gat));
  OR2_X1    g648(.A1(new_n814_), .A2(new_n815_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n651_), .A2(new_n531_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n614_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n621_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n317_), .A3(new_n429_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n317_), .B(new_n853_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(G169gat), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n856_), .A2(new_n858_), .A3(new_n861_), .ZN(G1348gat));
  NAND2_X1  g661(.A1(new_n806_), .A2(new_n620_), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n863_), .A2(new_n430_), .A3(new_n283_), .A4(new_n852_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n855_), .A2(new_n821_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n430_), .ZN(G1349gat));
  NOR2_X1   g665(.A1(new_n852_), .A2(new_n344_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n780_), .A2(new_n790_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n777_), .A2(KEYINPUT118), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n345_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n620_), .B(new_n867_), .C1(new_n870_), .C2(new_n815_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n806_), .A2(KEYINPUT123), .A3(new_n620_), .A4(new_n867_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n425_), .A3(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n344_), .A2(new_n491_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n853_), .B(new_n876_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n875_), .A2(KEYINPUT124), .A3(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1350gat));
  OAI21_X1  g681(.A(G190gat), .B1(new_n854_), .B2(new_n798_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n589_), .A2(new_n490_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n854_), .B2(new_n884_), .ZN(G1351gat));
  AND2_X1   g684(.A1(new_n837_), .A2(new_n851_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n317_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n821_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT125), .B(G204gat), .Z(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1353gat));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n345_), .B1(new_n892_), .B2(new_n327_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT126), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n886_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n892_), .A2(new_n327_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1354gat));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n886_), .B2(new_n583_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n837_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n851_), .ZN(new_n902_));
  NOR4_X1   g701(.A1(new_n901_), .A2(G218gat), .A3(new_n590_), .A4(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n898_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n886_), .A2(new_n899_), .A3(new_n589_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n901_), .A2(new_n798_), .A3(new_n902_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n905_), .B(KEYINPUT127), .C1(new_n899_), .C2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(G1355gat));
endmodule


