//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n839_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n207_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n213_), .B(new_n214_), .C1(new_n215_), .C2(KEYINPUT7), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n217_), .B(KEYINPUT66), .C1(G99gat), .C2(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT65), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n212_), .A2(new_n219_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  INV_X1    g023(.A(G92gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n216_), .A2(new_n218_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT8), .B1(new_n231_), .B2(new_n228_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(KEYINPUT64), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT64), .B1(new_n234_), .B2(new_n235_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n214_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n226_), .A2(KEYINPUT9), .A3(new_n227_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n227_), .A2(KEYINPUT9), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n239_), .A2(new_n222_), .A3(new_n212_), .A4(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n233_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G29gat), .B(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT69), .B(KEYINPUT15), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n220_), .A2(new_n221_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n219_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n228_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(KEYINPUT8), .A2(new_n255_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n212_), .A2(new_n222_), .A3(new_n241_), .A4(new_n240_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n234_), .A2(new_n235_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(G106gat), .B1(new_n260_), .B2(new_n236_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT67), .B1(new_n256_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n233_), .A2(new_n264_), .A3(new_n243_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n247_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n250_), .B(new_n251_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G232gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT34), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT35), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n272_), .B(new_n250_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n270_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n271_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT35), .B1(new_n271_), .B2(new_n274_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n206_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n272_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n271_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n205_), .B(KEYINPUT36), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT71), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n202_), .B1(new_n277_), .B2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n277_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n202_), .B2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT75), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G155gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G183gat), .B(G211gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT17), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G8gat), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G15gat), .B(G22gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G8gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n299_), .B(KEYINPUT73), .ZN(new_n304_));
  INV_X1    g103(.A(new_n302_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G57gat), .B(G64gat), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n308_), .A2(KEYINPUT11), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT11), .ZN(new_n310_));
  XOR2_X1   g109(.A(G71gat), .B(G78gat), .Z(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G231gat), .A2(G233gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n307_), .B(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n294_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(KEYINPUT17), .A3(new_n293_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n287_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT76), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n263_), .A2(new_n265_), .A3(new_n314_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n314_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n244_), .A2(KEYINPUT12), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n314_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n323_), .B(new_n325_), .C1(new_n326_), .C2(KEYINPUT12), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G230gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n256_), .A2(KEYINPUT67), .A3(new_n262_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n264_), .B1(new_n233_), .B2(new_n243_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n324_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n328_), .B1(new_n333_), .B2(new_n323_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G120gat), .B(G148gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT5), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G176gat), .B(G204gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT13), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n341_), .B(new_n342_), .C1(KEYINPUT68), .C2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G113gat), .B(G141gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT78), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G169gat), .B(G197gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  NAND2_X1  g151(.A1(G229gat), .A2(G233gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n303_), .A2(new_n306_), .A3(new_n247_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n247_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n354_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n307_), .A2(new_n249_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n353_), .A4(new_n355_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT77), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n352_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  AND4_X1   g164(.A1(new_n364_), .A2(new_n361_), .A3(new_n358_), .A4(new_n352_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n348_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT83), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G71gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(new_n213_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(KEYINPUT23), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n374_), .B(KEYINPUT81), .ZN(new_n377_));
  AOI211_X1 g176(.A(new_n373_), .B(new_n376_), .C1(new_n377_), .C2(KEYINPUT23), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT82), .B1(new_n380_), .B2(G169gat), .ZN(new_n381_));
  AOI21_X1  g180(.A(G176gat), .B1(new_n380_), .B2(G169gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n380_), .A2(KEYINPUT82), .A3(G169gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n379_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT26), .B(G190gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(G183gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT25), .B(G183gat), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n386_), .B(new_n389_), .C1(new_n390_), .C2(new_n387_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT24), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n393_));
  INV_X1    g192(.A(G169gat), .ZN(new_n394_));
  INV_X1    g193(.A(G176gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n392_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n396_), .A2(KEYINPUT24), .A3(new_n398_), .A4(new_n379_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n391_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT23), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n375_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n377_), .B2(new_n403_), .ZN(new_n405_));
  OAI22_X1  g204(.A1(new_n378_), .A2(new_n385_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n372_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G127gat), .B(G134gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G113gat), .B(G120gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n407_), .B(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n412_), .B(KEYINPUT84), .Z(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT30), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT31), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n411_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417_));
  INV_X1    g216(.A(G141gat), .ZN(new_n418_));
  INV_X1    g217(.A(G148gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G141gat), .A2(G148gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT2), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(KEYINPUT1), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT1), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(G155gat), .A3(G162gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n433_), .A3(new_n427_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n418_), .A2(new_n419_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n421_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT28), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G22gat), .B(G50gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G211gat), .B(G218gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(G197gat), .B(G204gat), .Z(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(KEYINPUT21), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G197gat), .B(G204gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT21), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n448_), .A2(KEYINPUT85), .A3(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n447_), .B(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n439_), .B2(new_n438_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(G228gat), .A3(G233gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G228gat), .A2(G233gat), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n451_), .B(new_n454_), .C1(new_n439_), .C2(new_n438_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n457_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(KEYINPUT86), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(KEYINPUT86), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n444_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n456_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n453_), .A2(new_n455_), .A3(KEYINPUT87), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n457_), .A3(new_n467_), .ZN(new_n468_));
  OR3_X1    g267(.A1(new_n456_), .A2(new_n463_), .A3(new_n457_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n464_), .A2(new_n443_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n462_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G1gat), .B(G29gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G85gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n410_), .A2(new_n436_), .A3(new_n430_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n408_), .A2(new_n409_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n408_), .A2(new_n409_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n437_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n482_), .A3(KEYINPUT91), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n438_), .A2(new_n484_), .A3(new_n410_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n485_), .A3(KEYINPUT4), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G225gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT92), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(KEYINPUT93), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n490_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n491_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n497_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(KEYINPUT93), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n477_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT98), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n498_), .A2(KEYINPUT93), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n494_), .B1(new_n498_), .B2(KEYINPUT93), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n476_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G226gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT19), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT89), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT20), .B1(new_n406_), .B2(new_n451_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n446_), .A2(new_n510_), .A3(KEYINPUT21), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n447_), .B(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n376_), .B1(new_n377_), .B2(KEYINPUT23), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n392_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n386_), .A2(new_n390_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n515_), .A2(KEYINPUT90), .A3(new_n401_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT90), .B1(new_n515_), .B2(new_n401_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n513_), .B(new_n514_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT22), .B(G169gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n395_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n379_), .B(new_n520_), .C1(new_n405_), .C2(new_n373_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n512_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n508_), .B1(new_n509_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n406_), .A2(new_n451_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n518_), .A2(new_n512_), .A3(new_n521_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n507_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(KEYINPUT20), .A4(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G8gat), .B(G36gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT18), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G64gat), .B(G92gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n533_), .A2(KEYINPUT32), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n509_), .A2(new_n522_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n508_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT97), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n525_), .A2(new_n539_), .A3(KEYINPUT20), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n539_), .B1(new_n525_), .B2(KEYINPUT20), .ZN(new_n541_));
  INV_X1    g340(.A(new_n524_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n538_), .B1(new_n543_), .B2(new_n526_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n535_), .B1(new_n544_), .B2(new_n534_), .ZN(new_n545_));
  OAI211_X1 g344(.A(KEYINPUT98), .B(new_n477_), .C1(new_n496_), .C2(new_n499_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n505_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n483_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n485_), .ZN(new_n549_));
  OR3_X1    g348(.A1(new_n548_), .A2(new_n549_), .A3(KEYINPUT95), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT95), .B1(new_n548_), .B2(new_n549_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n491_), .A3(new_n551_), .ZN(new_n552_));
  AOI211_X1 g351(.A(KEYINPUT96), .B(new_n493_), .C1(new_n486_), .C2(new_n488_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n552_), .B(new_n477_), .C1(new_n553_), .C2(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n523_), .A2(new_n533_), .A3(new_n527_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n533_), .B1(new_n523_), .B2(new_n527_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT33), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n504_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n504_), .A2(new_n561_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n547_), .A2(KEYINPUT99), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT99), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n505_), .A2(new_n545_), .A3(new_n566_), .A4(new_n546_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n471_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n505_), .A2(new_n546_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n525_), .A2(KEYINPUT20), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT97), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n525_), .A2(new_n539_), .A3(KEYINPUT20), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n572_), .A3(new_n524_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n573_), .A2(new_n507_), .B1(new_n537_), .B2(new_n536_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT100), .B1(new_n574_), .B2(new_n533_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT100), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n544_), .A2(new_n576_), .A3(new_n532_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT27), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n557_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT101), .B1(new_n559_), .B2(KEYINPUT27), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n582_), .B(new_n578_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  AND4_X1   g383(.A1(new_n569_), .A2(new_n471_), .A3(new_n580_), .A4(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n416_), .B1(new_n568_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n569_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n416_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n580_), .A2(new_n584_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n471_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n368_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n322_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n296_), .A3(new_n587_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT102), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT38), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n286_), .A2(new_n320_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT103), .Z(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n600_), .B2(new_n569_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n596_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n601_), .A3(new_n602_), .ZN(G1324gat));
  NAND3_X1  g402(.A1(new_n593_), .A2(new_n295_), .A3(new_n589_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT104), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n599_), .A2(new_n589_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(G8gat), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT39), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(KEYINPUT39), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n606_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n606_), .A2(new_n610_), .A3(KEYINPUT40), .A4(new_n609_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1325gat));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n416_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n593_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n599_), .B(KEYINPUT103), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n616_), .B1(new_n619_), .B2(new_n617_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n620_), .A2(new_n621_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n622_), .B2(new_n623_), .ZN(G1326gat));
  INV_X1    g423(.A(G22gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n593_), .A2(new_n625_), .A3(new_n471_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n471_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G22gat), .B1(new_n600_), .B2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n628_), .A2(KEYINPUT42), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(KEYINPUT42), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(G1327gat));
  NAND2_X1  g430(.A1(new_n277_), .A2(new_n285_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n320_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n592_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(G29gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n587_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n368_), .A2(new_n633_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n547_), .A2(KEYINPUT99), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n563_), .A2(new_n564_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n567_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n585_), .B1(new_n642_), .B2(new_n627_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n591_), .B1(new_n643_), .B2(new_n617_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n284_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT106), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n645_), .B(new_n646_), .C1(KEYINPUT37), .C2(new_n632_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n632_), .A2(KEYINPUT37), .ZN(new_n648_));
  OAI21_X1  g447(.A(KEYINPUT106), .B1(new_n648_), .B2(new_n284_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n639_), .B1(new_n644_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n287_), .A2(new_n639_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT44), .B(new_n638_), .C1(new_n651_), .C2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n638_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(KEYINPUT107), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT107), .B1(new_n655_), .B2(new_n656_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n587_), .B(new_n654_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT108), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(G29gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n660_), .B2(G29gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n637_), .B1(new_n662_), .B2(new_n663_), .ZN(G1328gat));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n654_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n655_), .A2(new_n656_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n667_), .B1(new_n670_), .B2(new_n657_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n666_), .B1(new_n671_), .B2(new_n589_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n635_), .A2(new_n666_), .A3(new_n589_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT45), .Z(new_n674_));
  OAI21_X1  g473(.A(new_n665_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n674_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n589_), .B(new_n654_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(new_n678_), .A3(KEYINPUT46), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(G1329gat));
  AND2_X1   g479(.A1(new_n617_), .A2(G43gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n671_), .A2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n635_), .A2(new_n617_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(G43gat), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT47), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n682_), .A2(new_n687_), .A3(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1330gat));
  AOI21_X1  g488(.A(G50gat), .B1(new_n635_), .B2(new_n471_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n471_), .A2(G50gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n671_), .B2(new_n691_), .ZN(G1331gat));
  NOR2_X1   g491(.A1(new_n348_), .A2(new_n367_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(new_n598_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G57gat), .B1(new_n697_), .B2(new_n569_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n348_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n322_), .A2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT109), .ZN(new_n701_));
  INV_X1    g500(.A(new_n367_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n644_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n569_), .A2(G57gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n698_), .B1(new_n703_), .B2(new_n704_), .ZN(G1332gat));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n696_), .B2(new_n589_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n589_), .A2(new_n706_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n703_), .B2(new_n710_), .ZN(G1333gat));
  INV_X1    g510(.A(G71gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n696_), .B2(new_n617_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT49), .Z(new_n714_));
  NAND2_X1  g513(.A1(new_n617_), .A2(new_n712_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n703_), .B2(new_n715_), .ZN(G1334gat));
  OAI21_X1  g515(.A(G78gat), .B1(new_n697_), .B2(new_n627_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT50), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n627_), .A2(G78gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n703_), .B2(new_n719_), .ZN(G1335gat));
  AND2_X1   g519(.A1(new_n695_), .A2(new_n634_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n224_), .A3(new_n587_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n694_), .A2(new_n633_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n587_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n722_), .B1(new_n727_), .B2(new_n224_), .ZN(G1336gat));
  INV_X1    g527(.A(new_n589_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G92gat), .B1(new_n724_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n721_), .A2(new_n225_), .A3(new_n589_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT111), .Z(G1337gat));
  OAI211_X1 g532(.A(new_n721_), .B(new_n617_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT112), .Z(new_n735_));
  OAI21_X1  g534(.A(G99gat), .B1(new_n724_), .B2(new_n416_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT51), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n736_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1338gat));
  OAI21_X1  g540(.A(G106gat), .B1(new_n724_), .B2(new_n627_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT52), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n721_), .A2(new_n214_), .A3(new_n471_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1339gat));
  NAND3_X1  g548(.A1(new_n321_), .A2(new_n702_), .A3(new_n348_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT54), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n341_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(new_n330_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n323_), .A2(new_n325_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT12), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n333_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n756_), .A2(new_n758_), .A3(KEYINPUT55), .A4(new_n328_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n339_), .B1(new_n755_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n756_), .A2(new_n758_), .A3(new_n328_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n328_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n753_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n759_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n339_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n752_), .B1(new_n763_), .B2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n362_), .A2(new_n364_), .A3(new_n352_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n353_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n352_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n359_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n770_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n342_), .B2(new_n341_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n632_), .B1(new_n769_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n778_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n339_), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n762_), .B(new_n340_), .C1(new_n766_), .C2(new_n759_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n761_), .A2(new_n785_), .A3(new_n762_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n775_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n341_), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n782_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n763_), .A2(KEYINPUT114), .A3(new_n768_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n775_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(KEYINPUT58), .A3(new_n792_), .A4(new_n787_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n287_), .A3(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n780_), .A2(new_n781_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n320_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n751_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n617_), .A2(new_n590_), .A3(new_n587_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(G113gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n367_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  INV_X1    g602(.A(new_n799_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n797_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n794_), .A2(new_n781_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n779_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n794_), .A2(KEYINPUT115), .A3(new_n781_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n806_), .B1(new_n811_), .B2(new_n633_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n633_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT116), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n751_), .A3(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n702_), .B(new_n805_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n802_), .B1(new_n817_), .B2(new_n801_), .ZN(G1340gat));
  INV_X1    g617(.A(G120gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n348_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n800_), .B(new_n820_), .C1(KEYINPUT60), .C2(new_n819_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n348_), .B(new_n805_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n819_), .ZN(G1341gat));
  AOI21_X1  g622(.A(G127gat), .B1(new_n800_), .B2(new_n633_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n805_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n633_), .A2(G127gat), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT117), .Z(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(new_n825_), .B2(new_n827_), .ZN(G1342gat));
  AOI21_X1  g627(.A(G134gat), .B1(new_n800_), .B2(new_n286_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n287_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT118), .B(G134gat), .Z(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n829_), .B1(new_n825_), .B2(new_n832_), .ZN(G1343gat));
  NAND4_X1  g632(.A1(new_n729_), .A2(new_n416_), .A3(new_n587_), .A4(new_n471_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT119), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n798_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n367_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n699_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n633_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT61), .B(G155gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1346gat));
  NOR3_X1   g642(.A1(new_n798_), .A2(new_n632_), .A3(new_n835_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(G162gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n650_), .A2(G162gat), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n798_), .A2(new_n835_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT120), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n847_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n849_), .B(new_n850_), .C1(G162gat), .C2(new_n844_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(G1347gat));
  NAND2_X1  g651(.A1(new_n588_), .A2(new_n589_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n471_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n751_), .B1(new_n813_), .B2(KEYINPUT116), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n806_), .B(new_n633_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n367_), .B(new_n854_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n394_), .B1(new_n858_), .B2(KEYINPUT62), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(KEYINPUT62), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n857_), .B(new_n859_), .C1(new_n858_), .C2(KEYINPUT62), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n815_), .A2(new_n367_), .A3(new_n519_), .A4(new_n854_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(G1348gat));
  NOR2_X1   g664(.A1(new_n798_), .A2(new_n471_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n853_), .A2(new_n395_), .A3(new_n348_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n699_), .B(new_n854_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n395_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(KEYINPUT122), .A3(new_n395_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n868_), .B1(new_n872_), .B2(new_n873_), .ZN(G1349gat));
  NOR2_X1   g673(.A1(new_n320_), .A2(new_n390_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n854_), .B(new_n875_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n876_), .A2(KEYINPUT123), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(KEYINPUT123), .ZN(new_n878_));
  NOR4_X1   g677(.A1(new_n798_), .A2(new_n471_), .A3(new_n320_), .A4(new_n853_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(G183gat), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n877_), .A2(new_n878_), .A3(new_n880_), .ZN(G1350gat));
  NAND2_X1  g680(.A1(new_n815_), .A2(new_n854_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G190gat), .B1(new_n882_), .B2(new_n830_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n286_), .A2(new_n386_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n882_), .B2(new_n884_), .ZN(G1351gat));
  NOR2_X1   g684(.A1(new_n627_), .A2(new_n587_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n416_), .A3(new_n589_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n797_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n367_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n348_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n894_), .A2(G204gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(G204gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n893_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n893_), .B2(new_n896_), .ZN(G1353gat));
  NAND3_X1  g697(.A1(new_n797_), .A2(new_n633_), .A3(new_n888_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT63), .B(G211gat), .Z(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT125), .B1(new_n899_), .B2(new_n901_), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n899_), .A2(KEYINPUT125), .A3(new_n901_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n899_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n899_), .A2(KEYINPUT126), .A3(new_n904_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n902_), .A2(new_n903_), .B1(new_n907_), .B2(new_n908_), .ZN(G1354gat));
  NOR3_X1   g708(.A1(new_n889_), .A2(G218gat), .A3(new_n632_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(G218gat), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n889_), .A2(new_n830_), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n911_), .B(KEYINPUT127), .C1(new_n912_), .C2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n912_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n910_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n914_), .A2(new_n917_), .ZN(G1355gat));
endmodule


