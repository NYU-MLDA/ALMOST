//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G106gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G85gat), .B(G92gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  INV_X1    g006(.A(G92gat), .ZN(new_n208_));
  OR3_X1    g007(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT9), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT6), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n206_), .A3(new_n209_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  OAI22_X1  g013(.A1(new_n214_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT65), .A3(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n211_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n205_), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n221_), .B(KEYINPUT66), .Z(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n219_), .B2(new_n205_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT67), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n213_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G29gat), .B(G36gat), .Z(new_n226_));
  XOR2_X1   g025(.A(G43gat), .B(G50gat), .Z(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT35), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G232gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT34), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n225_), .A2(new_n229_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n222_), .A2(new_n224_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n222_), .A2(KEYINPUT68), .A3(new_n224_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n213_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n228_), .B(KEYINPUT15), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n234_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n233_), .A2(new_n230_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI221_X1 g042(.A(new_n234_), .B1(new_n230_), .B2(new_n233_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G190gat), .B(G218gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G134gat), .B(G162gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT36), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT69), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n248_), .A2(KEYINPUT36), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n243_), .A2(new_n244_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n245_), .A2(new_n254_), .A3(new_n249_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n251_), .A2(new_n253_), .A3(new_n255_), .A4(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n253_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT37), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G1gat), .B(G8gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT72), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n264_), .A2(new_n265_), .ZN(new_n267_));
  INV_X1    g066(.A(G1gat), .ZN(new_n268_));
  INV_X1    g067(.A(G8gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT14), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n271_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G15gat), .B(G22gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  OR3_X1    g074(.A1(new_n266_), .A2(new_n267_), .A3(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n275_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n281_));
  XOR2_X1   g080(.A(G71gat), .B(G78gat), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n278_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT17), .ZN(new_n289_));
  XOR2_X1   g088(.A(G127gat), .B(G155gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G183gat), .B(G211gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n288_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT75), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n294_), .B(new_n289_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT76), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n288_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n261_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n283_), .A2(KEYINPUT12), .A3(new_n284_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n239_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n225_), .A2(new_n285_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n225_), .A2(new_n285_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(KEYINPUT12), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G230gat), .A2(G233gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n304_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(new_n305_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G120gat), .B(G148gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT5), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G176gat), .B(G204gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n309_), .A2(new_n312_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT13), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT13), .B1(new_n318_), .B2(new_n320_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n301_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT77), .Z(new_n327_));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n329_));
  INV_X1    g128(.A(G141gat), .ZN(new_n330_));
  INV_X1    g129(.A(G148gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G155gat), .B(G162gat), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n334_), .B(new_n335_), .C1(KEYINPUT1), .C2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(G141gat), .B2(G148gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n330_), .A2(new_n331_), .A3(KEYINPUT3), .ZN(new_n340_));
  AND3_X1   g139(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n339_), .A2(new_n340_), .B1(new_n341_), .B2(KEYINPUT86), .ZN(new_n342_));
  NAND3_X1  g141(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n343_), .A2(new_n344_), .B1(new_n333_), .B2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n336_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n337_), .B1(new_n347_), .B2(KEYINPUT87), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT87), .ZN(new_n349_));
  AOI211_X1 g148(.A(new_n349_), .B(new_n336_), .C1(new_n342_), .C2(new_n346_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n329_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n340_), .A2(new_n339_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n341_), .A2(KEYINPUT86), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n346_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n336_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n349_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n347_), .A2(KEYINPUT87), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT88), .A4(new_n337_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n351_), .A2(KEYINPUT29), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT93), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n362_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G197gat), .B(G204gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT21), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G197gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(G204gat), .ZN(new_n372_));
  INV_X1    g171(.A(G204gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G197gat), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n372_), .A2(new_n374_), .A3(KEYINPUT91), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT21), .B1(new_n372_), .B2(KEYINPUT91), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n370_), .B(new_n361_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n368_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(G228gat), .B2(G233gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n360_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n368_), .A2(KEYINPUT94), .A3(new_n377_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT94), .B1(new_n368_), .B2(new_n377_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n332_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n355_), .B2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n356_), .B2(new_n349_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n390_), .B2(new_n358_), .ZN(new_n391_));
  OAI211_X1 g190(.A(G228gat), .B(G233gat), .C1(new_n385_), .C2(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n381_), .A2(new_n382_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n382_), .B1(new_n381_), .B2(new_n392_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n328_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n381_), .A2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT95), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n381_), .A2(new_n392_), .A3(new_n382_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n328_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n400_), .A3(KEYINPUT90), .ZN(new_n401_));
  XOR2_X1   g200(.A(G22gat), .B(G50gat), .Z(new_n402_));
  NAND2_X1  g201(.A1(new_n351_), .A2(new_n359_), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n386_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n403_), .B2(new_n386_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n402_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n408_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n402_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n406_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n401_), .A2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n409_), .A2(new_n412_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(KEYINPUT90), .A3(new_n395_), .A4(new_n400_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n419_));
  OR2_X1    g218(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n420_));
  NAND2_X1  g219(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(G190gat), .A3(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT25), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G190gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT80), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G190gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n429_), .A3(KEYINPUT26), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT25), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G183gat), .ZN(new_n432_));
  AND4_X1   g231(.A1(new_n422_), .A2(new_n425_), .A3(new_n430_), .A4(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(KEYINPUT24), .A3(new_n435_), .ZN(new_n436_));
  OR3_X1    g235(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n437_));
  OR2_X1    g236(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n438_));
  NAND2_X1  g237(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n438_), .A2(new_n439_), .B1(G183gat), .B2(G190gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G183gat), .A2(G190gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(KEYINPUT23), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n436_), .B(new_n437_), .C1(new_n440_), .C2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n433_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(G169gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(KEYINPUT23), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT83), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n441_), .A2(new_n450_), .A3(KEYINPUT23), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n438_), .A2(new_n439_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n449_), .B(new_n451_), .C1(new_n452_), .C2(new_n441_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n423_), .A2(new_n427_), .A3(new_n429_), .A4(new_n424_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n447_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT84), .B1(new_n444_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n454_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n446_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n441_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n442_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n436_), .A2(new_n437_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n425_), .A2(new_n430_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n422_), .A2(new_n432_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n461_), .B(new_n462_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n458_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n456_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n419_), .B1(new_n468_), .B2(new_n378_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G226gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT19), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT25), .B(G183gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT26), .B(G190gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n436_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n453_), .A2(KEYINPUT96), .A3(new_n437_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT96), .B1(new_n453_), .B2(new_n437_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G183gat), .A2(G190gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n447_), .B1(new_n461_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n379_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT97), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT97), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n480_), .A2(new_n487_), .A3(new_n379_), .A4(new_n484_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n469_), .A2(new_n472_), .A3(new_n486_), .A4(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n453_), .A2(new_n437_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT96), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n453_), .A2(KEYINPUT96), .A3(new_n437_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n476_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n378_), .B1(new_n494_), .B2(new_n483_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n456_), .A2(new_n467_), .A3(new_n379_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(KEYINPUT20), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n471_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G8gat), .B(G36gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT18), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G64gat), .B(G92gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  AND3_X1   g301(.A1(new_n489_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n489_), .B2(new_n498_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n503_), .A2(new_n504_), .A3(KEYINPUT27), .ZN(new_n505_));
  INV_X1    g304(.A(new_n502_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n468_), .A2(new_n378_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n384_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n368_), .A2(new_n377_), .A3(KEYINPUT94), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n480_), .A2(new_n508_), .A3(new_n509_), .A4(new_n484_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(KEYINPUT20), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n471_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT20), .A4(new_n472_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT103), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n513_), .A2(KEYINPUT103), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n506_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT104), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n489_), .A2(new_n498_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n506_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n489_), .A2(new_n498_), .A3(KEYINPUT104), .A4(new_n502_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n505_), .B1(new_n522_), .B2(KEYINPUT27), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n418_), .A2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G127gat), .B(G134gat), .Z(new_n525_));
  XOR2_X1   g324(.A(G113gat), .B(G120gat), .Z(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT85), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  NAND3_X1  g328(.A1(new_n351_), .A2(new_n359_), .A3(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n525_), .A2(new_n526_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n390_), .B(new_n358_), .C1(new_n528_), .C2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(KEYINPUT4), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G225gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT4), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n351_), .A2(new_n536_), .A3(new_n359_), .A4(new_n529_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n530_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G29gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(G85gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT0), .B(G57gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n530_), .A2(KEYINPUT4), .A3(new_n532_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n537_), .A2(new_n535_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n539_), .B(new_n546_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G71gat), .B(G99gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(G43gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n468_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(new_n529_), .Z(new_n555_));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(G15gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT30), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT31), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n555_), .B(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n524_), .A2(new_n551_), .A3(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n523_), .A2(new_n417_), .A3(new_n550_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT100), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n537_), .A2(new_n534_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n547_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n530_), .A2(new_n532_), .A3(new_n535_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n544_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n564_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n533_), .A2(new_n534_), .A3(new_n537_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n570_), .A2(KEYINPUT100), .A3(new_n544_), .A4(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n503_), .A2(new_n504_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT33), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT99), .B1(new_n549_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n549_), .A2(KEYINPUT99), .A3(new_n575_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n544_), .A2(new_n575_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n539_), .B(new_n580_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT98), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n538_), .A2(new_n583_), .A3(new_n539_), .A4(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n574_), .A2(KEYINPUT101), .A3(new_n579_), .A4(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT101), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n572_), .A2(new_n585_), .A3(new_n573_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n549_), .A2(KEYINPUT99), .A3(new_n575_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n576_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n587_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n502_), .A2(KEYINPUT32), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n519_), .A2(KEYINPUT102), .A3(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT102), .B1(new_n519_), .B2(new_n592_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n593_), .A2(new_n550_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n586_), .A2(new_n591_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n563_), .B1(new_n597_), .B2(new_n417_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n562_), .B1(new_n598_), .B2(new_n561_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n278_), .B(new_n228_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n278_), .A2(new_n240_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n601_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n278_), .B2(new_n229_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n602_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G113gat), .B(G141gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G169gat), .B(G197gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n607_), .B(new_n608_), .Z(new_n609_));
  OR2_X1    g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n609_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT78), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n599_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n327_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n550_), .B(KEYINPUT105), .Z(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n268_), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n251_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n599_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n325_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n612_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n622_), .A2(new_n300_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G1gat), .B1(new_n625_), .B2(new_n551_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n619_), .A2(new_n626_), .ZN(new_n627_));
  MUX2_X1   g426(.A(new_n619_), .B(new_n627_), .S(KEYINPUT38), .Z(G1324gat));
  INV_X1    g427(.A(new_n523_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G8gat), .B1(new_n625_), .B2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(KEYINPUT106), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n327_), .A2(new_n269_), .A3(new_n523_), .A4(new_n615_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n630_), .A2(KEYINPUT106), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n631_), .A2(new_n636_), .A3(new_n632_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(G1325gat));
  INV_X1    g439(.A(new_n561_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G15gat), .B1(new_n625_), .B2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT41), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n616_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1326gat));
  INV_X1    g444(.A(G22gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n616_), .A2(new_n646_), .A3(new_n418_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G22gat), .B1(new_n625_), .B2(new_n417_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT108), .Z(G1327gat));
  INV_X1    g450(.A(new_n300_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n620_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n325_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n615_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G29gat), .B1(new_n655_), .B2(new_n550_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n325_), .A2(new_n300_), .A3(new_n612_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n599_), .A2(new_n659_), .A3(new_n261_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n599_), .B2(new_n261_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT44), .B(new_n658_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n618_), .A2(G29gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n656_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT111), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT112), .Z(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n655_), .A2(new_n674_), .A3(new_n523_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT45), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n629_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n599_), .A2(new_n261_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT43), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n599_), .A2(new_n261_), .A3(new_n659_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n657_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT109), .B1(new_n681_), .B2(KEYINPUT44), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n662_), .A2(new_n663_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT110), .B(new_n677_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT110), .B1(new_n664_), .B2(new_n677_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n673_), .B(new_n676_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n677_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(G36gat), .A3(new_n684_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n673_), .B1(new_n692_), .B2(new_n676_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n688_), .A2(new_n693_), .ZN(G1329gat));
  AND2_X1   g493(.A1(new_n561_), .A2(G43gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n664_), .A2(new_n667_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT113), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT113), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n664_), .A2(new_n698_), .A3(new_n667_), .A4(new_n695_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT114), .B(G43gat), .Z(new_n700_));
  INV_X1    g499(.A(new_n655_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n641_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n699_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT47), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n697_), .A2(new_n705_), .A3(new_n699_), .A4(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1330gat));
  AOI21_X1  g506(.A(G50gat), .B1(new_n655_), .B2(new_n418_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n418_), .A2(G50gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n668_), .B2(new_n709_), .ZN(G1331gat));
  NAND4_X1  g509(.A1(new_n621_), .A2(new_n652_), .A3(new_n622_), .A4(new_n613_), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n551_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT116), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n599_), .A2(new_n623_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n622_), .A3(new_n301_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT115), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n717_), .A2(new_n617_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n718_), .B2(new_n712_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n711_), .B2(new_n629_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT48), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n629_), .A2(G64gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n717_), .B2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n711_), .B2(new_n641_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n641_), .A2(G71gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n717_), .B2(new_n726_), .ZN(G1334gat));
  OAI21_X1  g526(.A(G78gat), .B1(new_n711_), .B2(new_n417_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT50), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n417_), .A2(G78gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n717_), .B2(new_n730_), .ZN(G1335gat));
  NAND2_X1  g530(.A1(new_n679_), .A2(new_n680_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n325_), .A2(new_n652_), .A3(new_n612_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n551_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n715_), .A2(new_n622_), .A3(new_n653_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n207_), .A3(new_n618_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1336gat));
  OAI21_X1  g537(.A(G92gat), .B1(new_n734_), .B2(new_n629_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n208_), .A3(new_n523_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n734_), .B2(new_n641_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n561_), .A2(new_n202_), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n742_), .A2(new_n743_), .B1(new_n736_), .B2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n745_), .B1(new_n743_), .B2(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n747_));
  OR2_X1    g546(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n746_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1338gat));
  XNOR2_X1  g550(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n752_));
  OAI21_X1  g551(.A(G106gat), .B1(new_n734_), .B2(new_n417_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT52), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT52), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n736_), .A2(new_n418_), .A3(new_n203_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n752_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n757_), .B(new_n752_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1339gat));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n301_), .A2(new_n762_), .A3(new_n325_), .A4(new_n613_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n325_), .A2(new_n613_), .A3(new_n652_), .A4(new_n260_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT54), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT57), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n612_), .A2(new_n320_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n310_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT55), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n309_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n307_), .A2(KEYINPUT55), .A3(new_n308_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n319_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n768_), .B1(new_n775_), .B2(KEYINPUT120), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT120), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n609_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n601_), .B1(new_n278_), .B2(new_n229_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n603_), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n606_), .B2(new_n609_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n776_), .A2(new_n778_), .B1(new_n321_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n620_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n767_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n771_), .A2(new_n772_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT120), .B(KEYINPUT56), .C1(new_n787_), .C2(new_n319_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n788_), .A2(new_n778_), .A3(new_n612_), .A4(new_n320_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n321_), .A2(new_n783_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT57), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n773_), .A2(new_n774_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n783_), .A2(new_n320_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n793_), .B1(new_n796_), .B2(new_n775_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n775_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n798_), .A2(KEYINPUT58), .A3(new_n794_), .A4(new_n795_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n797_), .A2(new_n799_), .A3(new_n261_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n786_), .A2(new_n792_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n766_), .B1(new_n801_), .B2(new_n300_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n524_), .A2(new_n618_), .A3(new_n561_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G113gat), .B1(new_n804_), .B2(new_n612_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n806_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n800_), .B1(new_n791_), .B2(KEYINPUT57), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n784_), .A2(new_n767_), .A3(new_n785_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n300_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n766_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n803_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(KEYINPUT59), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n810_), .A2(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n614_), .A2(G113gat), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n807_), .A2(new_n808_), .B1(new_n818_), .B2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n818_), .B2(new_n622_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n804_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n821_), .B1(new_n325_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(KEYINPUT60), .B2(new_n821_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT122), .B1(new_n822_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n325_), .B1(new_n810_), .B2(new_n817_), .ZN(new_n829_));
  OAI221_X1 g628(.A(new_n828_), .B1(new_n823_), .B2(new_n825_), .C1(new_n829_), .C2(new_n821_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(G1341gat));
  AOI21_X1  g630(.A(G127gat), .B1(new_n804_), .B2(new_n652_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n652_), .A2(G127gat), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT123), .Z(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n818_), .B2(new_n834_), .ZN(G1342gat));
  INV_X1    g634(.A(G134gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n804_), .A2(new_n836_), .A3(new_n785_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n260_), .B1(new_n810_), .B2(new_n817_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n836_), .ZN(G1343gat));
  NOR3_X1   g638(.A1(new_n617_), .A2(new_n417_), .A3(new_n523_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n815_), .A2(new_n641_), .A3(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n623_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(new_n330_), .ZN(G1344gat));
  NOR2_X1   g642(.A1(new_n841_), .A2(new_n325_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(new_n331_), .ZN(G1345gat));
  XNOR2_X1  g644(.A(KEYINPUT61), .B(G155gat), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT124), .B1(new_n841_), .B2(new_n300_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n841_), .A2(KEYINPUT124), .A3(new_n300_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n847_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n850_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n848_), .A3(new_n846_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1346gat));
  INV_X1    g653(.A(G162gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n841_), .A2(new_n855_), .A3(new_n260_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n841_), .A2(new_n620_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(G162gat), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT125), .B(new_n855_), .C1(new_n841_), .C2(new_n620_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n856_), .B1(new_n859_), .B2(new_n860_), .ZN(G1347gat));
  INV_X1    g660(.A(G169gat), .ZN(new_n862_));
  NOR4_X1   g661(.A1(new_n618_), .A2(new_n629_), .A3(new_n641_), .A4(new_n418_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n802_), .A2(new_n623_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n862_), .B1(new_n865_), .B2(KEYINPUT126), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n864_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT126), .B1(new_n868_), .B2(new_n612_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n866_), .A2(new_n867_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n866_), .B2(new_n870_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n868_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT22), .B(G169gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n612_), .A2(new_n874_), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT127), .Z(new_n876_));
  OAI22_X1  g675(.A1(new_n871_), .A2(new_n872_), .B1(new_n873_), .B2(new_n876_), .ZN(G1348gat));
  NAND2_X1  g676(.A1(new_n868_), .A2(new_n622_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g678(.A1(new_n423_), .A2(new_n424_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n868_), .A2(new_n652_), .ZN(new_n881_));
  MUX2_X1   g680(.A(new_n473_), .B(new_n880_), .S(new_n881_), .Z(G1350gat));
  OAI21_X1  g681(.A(G190gat), .B1(new_n873_), .B2(new_n260_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n868_), .A2(new_n474_), .A3(new_n785_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1351gat));
  NAND3_X1  g684(.A1(new_n418_), .A2(new_n551_), .A3(new_n523_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n802_), .A2(new_n561_), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n612_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n622_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g690(.A1(new_n887_), .A2(new_n652_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  AND2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n892_), .B2(new_n893_), .ZN(G1354gat));
  INV_X1    g695(.A(G218gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n887_), .A2(new_n897_), .A3(new_n785_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n887_), .A2(new_n261_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1355gat));
endmodule


