//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  INV_X1    g001(.A(G120gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G113gat), .ZN(new_n204_));
  INV_X1    g003(.A(G113gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G120gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G127gat), .B(G134gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(new_n204_), .A3(new_n206_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT31), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT80), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT25), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(G183gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT25), .B1(new_n217_), .B2(KEYINPUT80), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OR3_X1    g026(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n232_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(KEYINPUT82), .A3(new_n228_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n219_), .A2(KEYINPUT81), .A3(new_n224_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n227_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n220_), .A2(KEYINPUT22), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT22), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G169gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n245_), .A3(new_n221_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT83), .ZN(new_n247_));
  INV_X1    g046(.A(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n217_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n231_), .A2(new_n249_), .A3(new_n232_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n250_), .A3(new_n223_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n242_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G71gat), .B(G99gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G43gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n252_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(G15gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT30), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n255_), .B(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n212_), .B1(new_n259_), .B2(KEYINPUT84), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(KEYINPUT84), .B2(new_n259_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n259_), .A2(KEYINPUT84), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n212_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT27), .ZN(new_n265_));
  XOR2_X1   g064(.A(G8gat), .B(G36gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n248_), .A2(KEYINPUT26), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT26), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n217_), .A2(KEYINPUT25), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n215_), .A2(G183gat), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n271_), .A2(new_n273_), .A3(new_n274_), .A4(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n276_), .A2(new_n238_), .A3(new_n224_), .A4(new_n228_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT91), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n228_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n280_), .A2(KEYINPUT91), .A3(new_n224_), .A4(new_n276_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n223_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n283_), .B2(new_n221_), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT92), .B1(new_n284_), .B2(new_n250_), .ZN(new_n285_));
  AND4_X1   g084(.A1(KEYINPUT92), .A2(new_n250_), .A3(new_n223_), .A4(new_n246_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n279_), .B(new_n281_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G197gat), .B(G204gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G211gat), .B(G218gat), .ZN(new_n289_));
  OAI211_X1 g088(.A(KEYINPUT21), .B(new_n288_), .C1(new_n289_), .C2(KEYINPUT88), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291_));
  XOR2_X1   g090(.A(G211gat), .B(G218gat), .Z(new_n292_));
  INV_X1    g091(.A(KEYINPUT88), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G197gat), .B(G204gat), .Z(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(KEYINPUT21), .B2(new_n289_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n290_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n287_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n242_), .A2(new_n299_), .A3(new_n251_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n300_), .A3(KEYINPUT20), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT19), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n299_), .B1(new_n242_), .B2(new_n251_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n285_), .A2(new_n286_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n307_), .A2(new_n299_), .A3(new_n279_), .A4(new_n281_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT20), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n270_), .B1(new_n304_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n303_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n309_), .B1(new_n287_), .B2(new_n297_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n313_), .B1(new_n314_), .B2(new_n300_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n310_), .B1(new_n287_), .B2(new_n297_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(new_n305_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n270_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n265_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n270_), .B(KEYINPUT98), .Z(new_n321_));
  NOR2_X1   g120(.A1(new_n301_), .A2(new_n303_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n284_), .A2(new_n250_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT96), .B1(new_n323_), .B2(new_n277_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(new_n297_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n277_), .A3(KEYINPUT96), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n309_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n313_), .B1(new_n306_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n321_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n304_), .A2(new_n311_), .A3(new_n270_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(KEYINPUT27), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n320_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G155gat), .ZN(new_n336_));
  INV_X1    g135(.A(G162gat), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT85), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n343_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT2), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(G141gat), .A3(G148gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350_));
  NOR2_X1   g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n347_), .A2(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n340_), .B1(new_n345_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n351_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n346_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n339_), .B1(new_n338_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT1), .B1(new_n336_), .B2(new_n337_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n355_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G22gat), .B(G50gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n335_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n334_), .A3(new_n364_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT89), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n297_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n374_));
  AND2_X1   g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n297_), .B2(KEYINPUT87), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  OAI221_X1 g176(.A(new_n297_), .B1(KEYINPUT87), .B2(new_n375_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n373_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n378_), .A3(new_n373_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n370_), .A2(KEYINPUT90), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n377_), .A2(new_n378_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT90), .B1(new_n383_), .B2(new_n372_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n367_), .A2(new_n369_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n377_), .A2(new_n373_), .A3(new_n378_), .ZN(new_n386_));
  OAI22_X1  g185(.A1(new_n384_), .A2(new_n385_), .B1(new_n379_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n333_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n338_), .A2(new_n339_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n351_), .A2(new_n350_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n348_), .B1(G141gat), .B2(G148gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n346_), .A2(KEYINPUT2), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n342_), .A2(new_n344_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n391_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n356_), .A2(G155gat), .A3(G162gat), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n358_), .B(new_n398_), .C1(G155gat), .C2(G162gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n354_), .A3(new_n346_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n211_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n390_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n208_), .A2(new_n210_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n397_), .A2(new_n400_), .A3(new_n211_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT4), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n406_), .A3(new_n390_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G85gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(KEYINPUT0), .B(G57gat), .Z(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n412_), .B(new_n413_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n408_), .A2(new_n409_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n264_), .A2(new_n389_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n304_), .A2(new_n311_), .A3(new_n420_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n418_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n318_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT94), .B1(new_n330_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n397_), .A2(new_n400_), .A3(new_n211_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n429_), .A2(new_n401_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n407_), .A2(new_n403_), .B1(new_n430_), .B2(new_n390_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n428_), .B1(new_n431_), .B2(new_n416_), .ZN(new_n432_));
  AND4_X1   g231(.A1(new_n428_), .A2(new_n408_), .A3(new_n409_), .A4(new_n416_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n390_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n435_), .A2(new_n407_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT95), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n405_), .A2(new_n406_), .A3(new_n434_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n414_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n436_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n416_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n407_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT95), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI22_X1  g242(.A1(new_n432_), .A2(new_n433_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n427_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n330_), .A2(new_n426_), .A3(KEYINPUT94), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n425_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n382_), .A2(new_n387_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT97), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT94), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n417_), .A2(KEYINPUT33), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n431_), .A2(new_n428_), .A3(new_n416_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n437_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n441_), .A2(KEYINPUT95), .A3(new_n442_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n452_), .A2(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n446_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n448_), .B1(new_n457_), .B2(new_n424_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT97), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n388_), .A2(new_n418_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n333_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n449_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n419_), .B1(new_n463_), .B2(new_n264_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT10), .B(G99gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n467_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G85gat), .B(G92gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n471_), .A2(KEYINPUT66), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n474_), .A2(new_n477_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n465_), .B(KEYINPUT6), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(G106gat), .B2(new_n469_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n480_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n485_));
  OR3_X1    g284(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n475_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n492_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n479_), .B(new_n484_), .C1(new_n493_), .C2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G71gat), .B(G78gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n497_), .B1(KEYINPUT11), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT68), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n500_), .A3(KEYINPUT11), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n498_), .B2(KEYINPUT11), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n499_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT68), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n497_), .A4(new_n501_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT12), .B1(new_n496_), .B2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n496_), .A2(new_n510_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G230gat), .A2(G233gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(KEYINPUT64), .Z(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n481_), .A2(new_n483_), .A3(new_n480_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT66), .B1(new_n471_), .B2(new_n478_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT69), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n489_), .B(new_n492_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT69), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n484_), .A2(new_n479_), .A3(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT12), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n509_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n504_), .A2(new_n508_), .A3(KEYINPUT70), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n524_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n523_), .A2(new_n528_), .A3(KEYINPUT71), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT71), .B1(new_n523_), .B2(new_n528_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n513_), .B(new_n516_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n496_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(new_n509_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n515_), .B1(new_n533_), .B2(new_n512_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G120gat), .B(G148gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n535_), .A2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT13), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT13), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n542_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT76), .B(G8gat), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n551_), .B2(G1gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT77), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G15gat), .B(G22gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G1gat), .B(G8gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n556_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G29gat), .B(G36gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G43gat), .B(G50gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT79), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n559_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n559_), .A2(new_n563_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n556_), .B(new_n557_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n562_), .B(KEYINPUT15), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n568_), .A2(new_n571_), .A3(new_n565_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n567_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G169gat), .B(G197gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n567_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n549_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n464_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT35), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n532_), .A2(new_n562_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n523_), .A2(new_n570_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n586_), .A2(new_n583_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n587_), .B(new_n588_), .C1(new_n583_), .C2(new_n586_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT74), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT37), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n596_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n591_), .A2(new_n592_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n600_), .A3(KEYINPUT37), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(KEYINPUT70), .A3(KEYINPUT17), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(KEYINPUT17), .B2(new_n616_), .ZN(new_n618_));
  AND2_X1   g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n509_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n569_), .B(new_n620_), .ZN(new_n621_));
  MUX2_X1   g420(.A(new_n618_), .B(new_n617_), .S(new_n621_), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n610_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n582_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT99), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n582_), .A2(new_n627_), .A3(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n418_), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n629_), .A2(G1gat), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n464_), .A2(new_n606_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n581_), .A2(new_n623_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT100), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n637_), .B2(new_n630_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n631_), .A2(new_n632_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n633_), .A2(new_n638_), .A3(new_n639_), .ZN(G1324gat));
  NAND3_X1  g439(.A1(new_n634_), .A2(new_n332_), .A3(new_n635_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT101), .B1(new_n641_), .B2(G8gat), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n641_), .A2(G8gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n333_), .A2(new_n551_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n626_), .A2(new_n628_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n642_), .A2(new_n643_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n647_), .A2(new_n648_), .A3(new_n650_), .A4(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n646_), .A2(new_n645_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n650_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT40), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n652_), .A2(new_n656_), .A3(new_n658_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  OAI21_X1  g461(.A(G15gat), .B1(new_n637_), .B2(new_n264_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n629_), .A2(G15gat), .A3(new_n264_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1326gat));
  XNOR2_X1  g465(.A(new_n388_), .B(KEYINPUT104), .ZN(new_n667_));
  OAI21_X1  g466(.A(G22gat), .B1(new_n637_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT42), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n667_), .A2(G22gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n629_), .B2(new_n670_), .ZN(G1327gat));
  NOR2_X1   g470(.A1(new_n605_), .A2(new_n622_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n582_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G29gat), .B1(new_n673_), .B2(new_n418_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n581_), .A2(new_n622_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n462_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT97), .B(new_n448_), .C1(new_n424_), .C2(new_n457_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n264_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n419_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n680_), .A2(KEYINPUT105), .A3(new_n681_), .A4(new_n610_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n464_), .B2(new_n609_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n609_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT105), .B1(new_n685_), .B2(new_n681_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n675_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT106), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n687_), .A2(KEYINPUT106), .A3(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT44), .B(new_n675_), .C1(new_n684_), .C2(new_n686_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(G29gat), .A3(new_n418_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n674_), .B1(new_n692_), .B2(new_n694_), .ZN(G1328gat));
  XNOR2_X1  g494(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n693_), .A2(new_n332_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698_));
  INV_X1    g497(.A(new_n264_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n332_), .A2(new_n388_), .A3(new_n418_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n330_), .A2(new_n426_), .A3(KEYINPUT94), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n701_), .A2(new_n427_), .A3(new_n444_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n388_), .B1(new_n702_), .B2(new_n425_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n700_), .B1(new_n703_), .B2(KEYINPUT97), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n699_), .B1(new_n704_), .B2(new_n460_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n681_), .B(new_n610_), .C1(new_n705_), .C2(new_n419_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n683_), .A3(new_n682_), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n698_), .B(KEYINPUT44), .C1(new_n709_), .C2(new_n675_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n697_), .B1(new_n710_), .B2(new_n689_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G36gat), .ZN(new_n712_));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n673_), .A2(new_n713_), .A3(new_n332_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n696_), .B1(new_n712_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n696_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n716_), .B(new_n719_), .C1(new_n711_), .C2(G36gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1329gat));
  NAND3_X1  g520(.A1(new_n693_), .A2(G43gat), .A3(new_n699_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G43gat), .B1(new_n673_), .B2(new_n699_), .ZN(new_n724_));
  OR3_X1    g523(.A1(new_n723_), .A2(KEYINPUT47), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT47), .B1(new_n723_), .B2(new_n724_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1330gat));
  INV_X1    g526(.A(G50gat), .ZN(new_n728_));
  INV_X1    g527(.A(new_n667_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n673_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n448_), .B(new_n693_), .C1(new_n710_), .C2(new_n689_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n731_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT108), .B1(new_n731_), .B2(G50gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n732_), .B2(new_n733_), .ZN(G1331gat));
  INV_X1    g533(.A(new_n549_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n622_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n634_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(G57gat), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(new_n630_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n464_), .A2(new_n580_), .A3(new_n549_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n624_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(KEYINPUT109), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(KEYINPUT109), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n418_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n740_), .B1(new_n745_), .B2(new_n739_), .ZN(G1332gat));
  OAI21_X1  g545(.A(G64gat), .B1(new_n738_), .B2(new_n333_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT48), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n333_), .A2(G64gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n742_), .B2(new_n749_), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n738_), .B2(new_n264_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n264_), .A2(G71gat), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT110), .Z(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n742_), .B2(new_n754_), .ZN(G1334gat));
  OAI21_X1  g554(.A(G78gat), .B1(new_n738_), .B2(new_n667_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n667_), .A2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n742_), .B2(new_n758_), .ZN(G1335gat));
  NAND2_X1  g558(.A1(new_n741_), .A2(new_n672_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT111), .ZN(new_n761_));
  AOI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n418_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n580_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n735_), .A2(new_n623_), .A3(new_n763_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n709_), .A2(KEYINPUT112), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n709_), .A2(KEYINPUT112), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n418_), .A2(G85gat), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT113), .Z(new_n769_));
  AOI21_X1  g568(.A(new_n762_), .B1(new_n767_), .B2(new_n769_), .ZN(G1336gat));
  INV_X1    g569(.A(G92gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n761_), .A2(new_n771_), .A3(new_n332_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n767_), .A2(new_n332_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(new_n771_), .ZN(G1337gat));
  NAND3_X1  g573(.A1(new_n761_), .A2(new_n470_), .A3(new_n699_), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n264_), .B(new_n764_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n776_));
  INV_X1    g575(.A(G99gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT51), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n775_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1338gat));
  XNOR2_X1  g581(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n764_), .A2(new_n388_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n709_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(G106gat), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT52), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n761_), .A2(new_n468_), .A3(new_n448_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n783_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n786_), .A2(KEYINPUT52), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n785_), .B2(G106gat), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n788_), .B(new_n783_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n789_), .A2(new_n794_), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n580_), .A2(new_n546_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n531_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT55), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n531_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n513_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n515_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n799_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n541_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n541_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n796_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n564_), .A2(new_n565_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n568_), .A2(new_n571_), .A3(new_n566_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n577_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n579_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n546_), .B2(new_n542_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n605_), .B1(new_n809_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n813_), .A2(new_n544_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n541_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n541_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n609_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT58), .B(new_n818_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT57), .B(new_n605_), .C1(new_n809_), .C2(new_n814_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n817_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n623_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n736_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n609_), .B1(new_n829_), .B2(KEYINPUT115), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831_));
  AOI211_X1 g630(.A(new_n831_), .B(new_n736_), .C1(new_n545_), .C2(new_n548_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT54), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n549_), .A2(new_n737_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n831_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n829_), .A2(KEYINPUT115), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n609_), .A4(new_n837_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n833_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n828_), .A2(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n264_), .A2(new_n389_), .A3(new_n630_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n205_), .A3(new_n580_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(KEYINPUT59), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n763_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n849_), .B2(new_n205_), .ZN(G1340gat));
  OAI21_X1  g649(.A(new_n203_), .B1(new_n549_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n844_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n203_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n549_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n203_), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n844_), .A2(new_n855_), .A3(new_n622_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n623_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n855_), .ZN(G1342gat));
  INV_X1    g657(.A(G134gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n843_), .B2(new_n605_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n861_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n846_), .A2(new_n848_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n609_), .A2(new_n859_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n862_), .A2(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1343gat));
  NOR3_X1   g665(.A1(new_n332_), .A2(new_n388_), .A3(new_n630_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n841_), .A2(new_n264_), .A3(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n763_), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n869_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n549_), .ZN(new_n871_));
  XOR2_X1   g670(.A(new_n871_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g671(.A1(new_n868_), .A2(new_n623_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT61), .B(G155gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n868_), .B2(new_n609_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n606_), .A2(new_n337_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n868_), .B2(new_n877_), .ZN(G1347gat));
  NAND3_X1  g677(.A1(new_n699_), .A2(new_n332_), .A3(new_n630_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n729_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n841_), .A2(new_n580_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(G169gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(G169gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(KEYINPUT118), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886_));
  AOI211_X1 g685(.A(new_n886_), .B(new_n882_), .C1(new_n881_), .C2(G169gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n841_), .A2(new_n880_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n580_), .A2(new_n283_), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT119), .Z(new_n890_));
  OAI22_X1  g689(.A1(new_n885_), .A2(new_n887_), .B1(new_n888_), .B2(new_n890_), .ZN(G1348gat));
  NAND2_X1  g690(.A1(new_n841_), .A2(new_n388_), .ZN(new_n892_));
  NOR4_X1   g691(.A1(new_n892_), .A2(new_n221_), .A3(new_n549_), .A4(new_n879_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n221_), .B1(new_n888_), .B2(new_n549_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n894_), .A2(KEYINPUT120), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(KEYINPUT120), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n895_), .B2(new_n896_), .ZN(G1349gat));
  OR3_X1    g696(.A1(new_n892_), .A2(new_n623_), .A3(new_n879_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n888_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n623_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n898_), .A2(new_n217_), .B1(new_n899_), .B2(new_n900_), .ZN(G1350gat));
  OAI21_X1  g700(.A(G190gat), .B1(new_n888_), .B2(new_n609_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n606_), .A2(new_n213_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n888_), .B2(new_n903_), .ZN(G1351gat));
  NAND2_X1  g703(.A1(new_n264_), .A2(new_n461_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n906_), .A2(KEYINPUT121), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(KEYINPUT121), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n332_), .A3(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n828_), .B2(new_n840_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n580_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n735_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g713(.A(new_n910_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n622_), .A2(new_n916_), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT122), .Z(new_n918_));
  NOR2_X1   g717(.A1(new_n915_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(KEYINPUT124), .B1(new_n919_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n923_), .B(new_n920_), .C1(new_n915_), .C2(new_n918_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n918_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n910_), .A2(new_n921_), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n927_), .ZN(new_n929_));
  AOI22_X1  g728(.A1(new_n922_), .A2(new_n924_), .B1(new_n928_), .B2(new_n929_), .ZN(G1354gat));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT126), .B(G218gat), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n909_), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n816_), .A2(new_n815_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n622_), .B1(new_n935_), .B2(new_n826_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n606_), .B(new_n934_), .C1(new_n936_), .C2(new_n839_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(KEYINPUT125), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n910_), .A2(new_n939_), .A3(new_n606_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n933_), .B1(new_n938_), .B2(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n910_), .A2(new_n610_), .A3(new_n933_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n931_), .B1(new_n941_), .B2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n939_), .B1(new_n910_), .B2(new_n606_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n839_), .B1(new_n827_), .B2(new_n623_), .ZN(new_n946_));
  NOR4_X1   g745(.A1(new_n946_), .A2(KEYINPUT125), .A3(new_n605_), .A4(new_n909_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n932_), .B1(new_n945_), .B2(new_n947_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n948_), .A2(KEYINPUT127), .A3(new_n942_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n944_), .A2(new_n949_), .ZN(G1355gat));
endmodule


