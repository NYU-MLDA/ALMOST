//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT90), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(KEYINPUT90), .A3(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  INV_X1    g011(.A(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n203_), .B1(new_n211_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT88), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT85), .A3(G183gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(KEYINPUT87), .A3(G190gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(G190gat), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n224_), .B(new_n226_), .C1(new_n227_), .C2(KEYINPUT86), .ZN(new_n228_));
  NAND2_X1  g027(.A1(KEYINPUT87), .A2(G190gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT86), .A3(KEYINPUT26), .ZN(new_n230_));
  NAND2_X1  g029(.A1(KEYINPUT85), .A2(G183gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT25), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n217_), .B(new_n222_), .C1(new_n228_), .C2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT89), .ZN(new_n235_));
  OR3_X1    g034(.A1(new_n204_), .A2(KEYINPUT89), .A3(KEYINPUT23), .ZN(new_n236_));
  OR3_X1    g035(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(KEYINPUT86), .A2(KEYINPUT26), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n240_), .A2(new_n229_), .B1(new_n231_), .B2(KEYINPUT25), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n213_), .A2(KEYINPUT26), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n241_), .A2(new_n224_), .A3(new_n226_), .A4(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n217_), .B1(new_n245_), .B2(new_n222_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n216_), .B1(new_n239_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT91), .B(KEYINPUT30), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n216_), .B(new_n248_), .C1(new_n239_), .C2(new_n246_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT92), .B(G43gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT94), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G134gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G127gat), .ZN(new_n259_));
  INV_X1    g058(.A(G127gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(G134gat), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n259_), .A2(new_n261_), .A3(KEYINPUT95), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT95), .B1(new_n259_), .B2(new_n261_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n257_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n261_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT95), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n259_), .A2(new_n261_), .A3(KEYINPUT95), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n256_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n254_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n250_), .A2(new_n271_), .A3(new_n251_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n255_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n270_), .B1(new_n255_), .B2(new_n272_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT31), .ZN(new_n276_));
  XOR2_X1   g075(.A(G71gat), .B(G99gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT93), .ZN(new_n278_));
  INV_X1    g077(.A(G15gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(G227gat), .A3(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n278_), .B(G15gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n276_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n281_), .A2(new_n276_), .A3(new_n284_), .ZN(new_n286_));
  OAI22_X1  g085(.A1(new_n274_), .A2(new_n275_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n275_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n286_), .A2(new_n285_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n273_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT99), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT99), .ZN(new_n295_));
  INV_X1    g094(.A(G204gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(G197gat), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n297_), .A2(KEYINPUT21), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G218gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G211gat), .ZN(new_n301_));
  INV_X1    g100(.A(G211gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G218gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT21), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(new_n293_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n293_), .A2(new_n305_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n299_), .A2(new_n306_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n216_), .B(new_n308_), .C1(new_n239_), .C2(new_n246_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n209_), .A2(new_n210_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n222_), .A2(new_n237_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n225_), .A2(G190gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n212_), .A2(KEYINPUT25), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n223_), .A2(G183gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n312_), .A2(new_n242_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT101), .A4(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT101), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n222_), .A3(new_n237_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(new_n211_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n235_), .A2(new_n236_), .A3(new_n214_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n316_), .A2(new_n319_), .B1(new_n203_), .B2(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n309_), .B(KEYINPUT20), .C1(new_n321_), .C2(new_n308_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT19), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G8gat), .B(G36gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT18), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G64gat), .B(G92gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n324_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT20), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n321_), .B2(new_n308_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n308_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n247_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n325_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT27), .ZN(new_n337_));
  INV_X1    g136(.A(new_n329_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT104), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT20), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n320_), .A2(new_n203_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n315_), .A2(new_n222_), .A3(new_n237_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT101), .B1(new_n343_), .B2(new_n310_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n318_), .A2(new_n211_), .A3(new_n317_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n342_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n341_), .B1(new_n346_), .B2(new_n333_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n347_), .A2(KEYINPUT104), .A3(new_n330_), .A4(new_n309_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n308_), .B(new_n342_), .C1(new_n211_), .C2(new_n318_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n334_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n324_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n340_), .A2(new_n348_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n337_), .B1(new_n338_), .B2(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(KEYINPUT97), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT97), .ZN(new_n358_));
  AND2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT96), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT96), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G141gat), .A3(G148gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G141gat), .ZN(new_n369_));
  INV_X1    g168(.A(G148gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT3), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n363_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT2), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n368_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n362_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n369_), .A2(new_n370_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n364_), .A2(new_n366_), .A3(new_n379_), .A4(new_n380_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n359_), .A2(new_n360_), .A3(KEYINPUT1), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT29), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n333_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n378_), .B2(new_n384_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n391_), .B2(new_n308_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n388_), .A2(new_n392_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n385_), .A2(KEYINPUT29), .ZN(new_n399_));
  XOR2_X1   g198(.A(KEYINPUT98), .B(KEYINPUT28), .Z(new_n400_));
  XNOR2_X1  g199(.A(G22gat), .B(G50gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n399_), .B(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n396_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(KEYINPUT100), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n398_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n357_), .A2(new_n361_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n371_), .A2(new_n373_), .B1(new_n375_), .B2(KEYINPUT2), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n368_), .B2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n269_), .B(new_n264_), .C1(new_n409_), .C2(new_n383_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n270_), .A2(new_n384_), .A3(new_n378_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(KEYINPUT4), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n270_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n385_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n412_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n410_), .A2(new_n413_), .A3(new_n411_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT102), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT102), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n410_), .A2(new_n411_), .A3(new_n421_), .A4(new_n413_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n418_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G85gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT0), .B(G57gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n425_), .B(new_n426_), .Z(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n418_), .A2(new_n420_), .A3(new_n427_), .A4(new_n422_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n395_), .A2(new_n403_), .A3(KEYINPUT100), .A4(new_n397_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n406_), .A2(new_n429_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT105), .B(KEYINPUT27), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n325_), .A2(new_n335_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n338_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n434_), .B1(new_n436_), .B2(new_n336_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n354_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n406_), .A2(new_n431_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n329_), .A2(KEYINPUT32), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n353_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n429_), .A2(new_n430_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n325_), .A2(new_n440_), .A3(new_n335_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n412_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n410_), .A2(new_n414_), .A3(new_n411_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n428_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT33), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n430_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n420_), .A2(new_n422_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n451_), .A2(KEYINPUT33), .A3(new_n427_), .A4(new_n418_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n450_), .A2(new_n452_), .A3(new_n336_), .A4(new_n436_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n439_), .B1(new_n445_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n292_), .B1(new_n438_), .B2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n354_), .A2(new_n437_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n443_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n406_), .A2(new_n431_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .A4(new_n291_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT76), .B(G8gat), .Z(new_n462_));
  INV_X1    g261(.A(G1gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G1gat), .B(G8gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n466_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G29gat), .B(G36gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G43gat), .B(G50gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT80), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n469_), .B(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(G229gat), .A3(G233gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n469_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n472_), .B(KEYINPUT15), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n469_), .A2(new_n474_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT81), .Z(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n461_), .B1(new_n476_), .B2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G113gat), .B(G141gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT82), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT83), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G169gat), .B(G197gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  AOI211_X1 g290(.A(new_n461_), .B(new_n491_), .C1(new_n476_), .C2(new_n483_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n460_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G190gat), .B(G218gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT75), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G134gat), .B(G162gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT36), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G232gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT74), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT6), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(G99gat), .A3(G106gat), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G85gat), .ZN(new_n512_));
  INV_X1    g311(.A(G92gat), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT9), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  INV_X1    g315(.A(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G85gat), .B(G92gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT9), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n515_), .A2(new_n518_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n508_), .A2(new_n510_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n519_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT8), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT65), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532_));
  INV_X1    g331(.A(G99gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n517_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n524_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n520_), .B1(new_n511_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT65), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT8), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n530_), .B(new_n520_), .C1(new_n511_), .C2(new_n535_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT64), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n527_), .A2(new_n528_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT64), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n530_), .A4(new_n520_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n523_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n472_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n531_), .A2(new_n538_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n522_), .A2(KEYINPUT68), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n515_), .A2(new_n550_), .A3(new_n518_), .A4(new_n521_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n478_), .B1(new_n548_), .B2(new_n552_), .ZN(new_n553_));
  AOI211_X1 g352(.A(new_n502_), .B(new_n506_), .C1(new_n547_), .C2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n506_), .A2(new_n502_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n547_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n506_), .A2(new_n502_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n501_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(new_n558_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n499_), .A2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n561_), .A2(new_n554_), .A3(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT37), .B1(new_n560_), .B2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n555_), .A2(new_n562_), .A3(new_n499_), .A4(new_n559_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n500_), .B1(new_n561_), .B2(new_n554_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G57gat), .B(G64gat), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT66), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G57gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(G64gat), .ZN(new_n575_));
  INV_X1    g374(.A(G64gat), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(G57gat), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n575_), .A2(new_n577_), .A3(KEYINPUT66), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT11), .B1(new_n573_), .B2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(new_n572_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT66), .B1(new_n575_), .B2(new_n577_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT11), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n579_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(KEYINPUT11), .B(new_n580_), .C1(new_n573_), .C2(new_n578_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT77), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n588_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n469_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G127gat), .B(G155gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT17), .Z(new_n598_));
  OR2_X1    g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(KEYINPUT17), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n592_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n570_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT79), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n495_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT67), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n546_), .B2(new_n588_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n546_), .A2(new_n588_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n588_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n610_), .B(KEYINPUT67), .C1(new_n548_), .C2(new_n523_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n546_), .B2(new_n588_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n610_), .B(KEYINPUT12), .C1(new_n548_), .C2(new_n552_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n613_), .A4(new_n609_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT5), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n615_), .A2(new_n619_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT71), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n615_), .A2(KEYINPUT71), .A3(new_n619_), .A4(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n623_), .B(KEYINPUT70), .Z(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT13), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(KEYINPUT13), .A3(new_n631_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(KEYINPUT72), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT72), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT13), .B1(new_n628_), .B2(new_n631_), .ZN(new_n638_));
  AOI211_X1 g437(.A(new_n633_), .B(new_n630_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n606_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n463_), .A3(new_n443_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT38), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n634_), .A2(new_n635_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n494_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n455_), .A2(new_n459_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n566_), .A2(new_n568_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .A4(new_n602_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT106), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n443_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n647_), .B1(new_n654_), .B2(G1gat), .ZN(new_n655_));
  AOI211_X1 g454(.A(KEYINPUT107), .B(new_n463_), .C1(new_n653_), .C2(new_n443_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n646_), .B1(new_n655_), .B2(new_n656_), .ZN(G1324gat));
  INV_X1    g456(.A(new_n456_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n462_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n643_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(KEYINPUT108), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n643_), .A2(new_n662_), .A3(new_n659_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n652_), .A2(new_n456_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(G8gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n664_), .B2(G8gat), .ZN(new_n667_));
  OAI22_X1  g466(.A1(new_n661_), .A2(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI221_X1 g469(.A(KEYINPUT40), .B1(new_n666_), .B2(new_n667_), .C1(new_n661_), .C2(new_n663_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  NAND3_X1  g471(.A1(new_n644_), .A2(new_n279_), .A3(new_n291_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n653_), .A2(new_n291_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n674_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT41), .B1(new_n674_), .B2(G15gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(G1326gat));
  OR3_X1    g476(.A1(new_n643_), .A2(G22gat), .A3(new_n458_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n653_), .A2(new_n439_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(G22gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G22gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(G1327gat));
  NOR3_X1   g482(.A1(new_n648_), .A2(new_n602_), .A3(new_n494_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(new_n570_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n650_), .B2(new_n686_), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT43), .B(new_n570_), .C1(new_n455_), .C2(new_n459_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT44), .B(new_n684_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n691_), .A2(G29gat), .A3(new_n443_), .A4(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(G29gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n651_), .A2(new_n602_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n648_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n495_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n698_), .B2(new_n457_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n693_), .A2(new_n699_), .ZN(G1328gat));
  NOR2_X1   g499(.A1(new_n456_), .A2(G36gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n495_), .A2(new_n697_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT110), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n495_), .A2(new_n704_), .A3(new_n697_), .A4(new_n701_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n703_), .A2(KEYINPUT45), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT45), .B1(new_n703_), .B2(new_n705_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n691_), .A2(new_n658_), .A3(new_n692_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G36gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G36gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT46), .B(new_n708_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  XNOR2_X1  g516(.A(KEYINPUT111), .B(G43gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n698_), .B2(new_n292_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n691_), .A2(new_n692_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n291_), .A2(G43gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n720_), .B2(new_n458_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n458_), .A2(G50gat), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT112), .Z(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n698_), .B2(new_n726_), .ZN(G1331gat));
  INV_X1    g526(.A(new_n602_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n493_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n650_), .A2(new_n651_), .A3(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(new_n641_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n457_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n493_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n605_), .A2(new_n648_), .A3(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n574_), .A3(new_n443_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(G1332gat));
  AOI21_X1  g536(.A(new_n576_), .B1(new_n731_), .B2(new_n658_), .ZN(new_n738_));
  XOR2_X1   g537(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n576_), .A3(new_n658_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n731_), .B2(new_n291_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT49), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n735_), .A2(new_n743_), .A3(new_n291_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1334gat));
  INV_X1    g546(.A(G78gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n735_), .A2(new_n748_), .A3(new_n439_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n731_), .A2(new_n439_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(G78gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT50), .B(new_n748_), .C1(new_n731_), .C2(new_n439_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT114), .ZN(G1335gat));
  NAND3_X1  g554(.A1(new_n648_), .A2(new_n728_), .A3(new_n494_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT43), .B1(new_n460_), .B2(new_n570_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n650_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n457_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT72), .B1(new_n634_), .B2(new_n635_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n638_), .A2(new_n639_), .A3(new_n637_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n695_), .B(new_n734_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n696_), .B1(new_n636_), .B2(new_n640_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT115), .A3(new_n734_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n512_), .A3(new_n443_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n761_), .A2(new_n770_), .ZN(G1336gat));
  OAI21_X1  g570(.A(G92gat), .B1(new_n760_), .B2(new_n456_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n513_), .A3(new_n658_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1337gat));
  AOI21_X1  g573(.A(new_n533_), .B1(new_n759_), .B2(new_n291_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n777_));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n291_), .A2(new_n516_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n778_), .B1(new_n769_), .B2(new_n780_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT116), .B(new_n779_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n776_), .B(new_n777_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(KEYINPUT118), .ZN(new_n784_));
  AND4_X1   g583(.A1(KEYINPUT115), .A2(new_n641_), .A3(new_n695_), .A4(new_n734_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT115), .B1(new_n767_), .B2(new_n734_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n780_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT116), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n769_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n775_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n790_), .B2(new_n777_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n784_), .B1(new_n792_), .B2(new_n794_), .ZN(G1338gat));
  NOR2_X1   g594(.A1(new_n638_), .A2(new_n639_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n796_), .A2(new_n602_), .A3(new_n493_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n439_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT119), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(G106gat), .B1(new_n798_), .B2(KEYINPUT119), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT52), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n759_), .A2(new_n803_), .A3(new_n439_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n804_), .A2(new_n799_), .A3(new_n805_), .A4(G106gat), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n802_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n769_), .A2(new_n517_), .A3(new_n439_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT53), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n811_), .A3(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n491_), .B1(new_n476_), .B2(new_n483_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n475_), .A2(new_n482_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n482_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n479_), .A2(new_n480_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n489_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n618_), .A2(new_n609_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n616_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n539_), .A2(new_n545_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n522_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n825_), .B2(new_n610_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n614_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n822_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n830_), .A2(KEYINPUT55), .A3(new_n613_), .A4(new_n617_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n619_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT121), .B(new_n614_), .C1(new_n822_), .C2(new_n826_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n829_), .A2(new_n831_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n629_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n835_), .A2(KEYINPUT56), .A3(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n628_), .A2(new_n493_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n821_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n651_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n814_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n820_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n835_), .A2(KEYINPUT56), .A3(new_n836_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT56), .B1(new_n835_), .B2(new_n836_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n570_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n841_), .A2(KEYINPUT58), .A3(new_n847_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n842_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT57), .B(new_n651_), .C1(new_n855_), .C2(new_n821_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n846_), .A2(new_n854_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n728_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n634_), .A2(new_n635_), .A3(new_n729_), .A4(new_n570_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n862_), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n658_), .A2(new_n292_), .A3(new_n457_), .A4(new_n439_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(G113gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n493_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n863_), .A2(KEYINPUT59), .A3(new_n864_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n494_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n872_), .B2(new_n867_), .ZN(G1340gat));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n796_), .B2(KEYINPUT60), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n866_), .B(new_n875_), .C1(KEYINPUT60), .C2(new_n874_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n642_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n874_), .ZN(G1341gat));
  NAND3_X1  g677(.A1(new_n866_), .A2(new_n260_), .A3(new_n602_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n728_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n260_), .ZN(G1342gat));
  XNOR2_X1  g680(.A(KEYINPUT123), .B(G134gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n686_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n258_), .B1(new_n865_), .B2(new_n651_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT122), .B(new_n258_), .C1(new_n865_), .C2(new_n651_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n884_), .B1(new_n887_), .B2(new_n888_), .ZN(G1343gat));
  AOI21_X1  g688(.A(new_n861_), .B1(new_n857_), .B2(new_n728_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n291_), .A2(new_n458_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n658_), .A2(new_n457_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(new_n493_), .A3(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n641_), .A3(new_n894_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g697(.A1(new_n893_), .A2(new_n602_), .A3(new_n894_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1346gat));
  NAND2_X1  g700(.A1(new_n893_), .A2(new_n894_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G162gat), .B1(new_n902_), .B2(new_n570_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n651_), .A2(G162gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n902_), .B2(new_n904_), .ZN(G1347gat));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n291_), .A2(new_n457_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n907_), .A2(new_n456_), .A3(new_n439_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n890_), .B2(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n651_), .B1(new_n855_), .B2(new_n821_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n911_), .A2(new_n814_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n602_), .B1(new_n912_), .B2(new_n856_), .ZN(new_n913_));
  OAI211_X1 g712(.A(KEYINPUT124), .B(new_n908_), .C1(new_n913_), .C2(new_n861_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n914_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT22), .B(G169gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n493_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n890_), .A2(new_n909_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n493_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n920_), .B2(G169gat), .ZN(new_n921_));
  AOI211_X1 g720(.A(KEYINPUT62), .B(new_n218_), .C1(new_n919_), .C2(new_n493_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n917_), .B1(new_n921_), .B2(new_n922_), .ZN(G1348gat));
  NOR2_X1   g722(.A1(new_n796_), .A2(G176gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n915_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n863_), .A2(new_n908_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G176gat), .B1(new_n926_), .B2(new_n642_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(KEYINPUT125), .A3(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929_));
  INV_X1    g728(.A(new_n924_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n910_), .B2(new_n914_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n219_), .B1(new_n919_), .B2(new_n641_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n929_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n928_), .A2(new_n933_), .ZN(G1349gat));
  AND2_X1   g733(.A1(new_n313_), .A2(new_n314_), .ZN(new_n935_));
  AOI211_X1 g734(.A(new_n935_), .B(new_n728_), .C1(new_n910_), .C2(new_n914_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n926_), .A2(new_n728_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G183gat), .B1(new_n937_), .B2(KEYINPUT126), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n939_), .B1(new_n926_), .B2(new_n728_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n936_), .B1(new_n938_), .B2(new_n940_), .ZN(G1350gat));
  INV_X1    g740(.A(new_n915_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n845_), .A2(new_n312_), .A3(new_n242_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n570_), .B1(new_n910_), .B2(new_n914_), .ZN(new_n944_));
  OAI22_X1  g743(.A1(new_n942_), .A2(new_n943_), .B1(new_n944_), .B2(new_n213_), .ZN(G1351gat));
  NOR2_X1   g744(.A1(new_n456_), .A2(new_n443_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n893_), .A2(new_n493_), .A3(new_n946_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n863_), .A2(new_n891_), .A3(new_n946_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n642_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(new_n296_), .ZN(G1353gat));
  XNOR2_X1  g750(.A(KEYINPUT63), .B(G211gat), .ZN(new_n952_));
  OR2_X1    g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n893_), .A2(new_n602_), .A3(new_n946_), .ZN(new_n954_));
  MUX2_X1   g753(.A(new_n952_), .B(new_n953_), .S(new_n954_), .Z(G1354gat));
  INV_X1    g754(.A(new_n946_), .ZN(new_n956_));
  NOR4_X1   g755(.A1(new_n890_), .A2(new_n570_), .A3(new_n892_), .A4(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n845_), .A2(new_n300_), .ZN(new_n958_));
  OAI22_X1  g757(.A1(new_n957_), .A2(new_n300_), .B1(new_n949_), .B2(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  OAI221_X1 g760(.A(KEYINPUT127), .B1(new_n949_), .B2(new_n958_), .C1(new_n957_), .C2(new_n300_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1355gat));
endmodule


