//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT29), .ZN(new_n204_));
  INV_X1    g003(.A(G155gat), .ZN(new_n205_));
  INV_X1    g004(.A(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G141gat), .ZN(new_n210_));
  INV_X1    g009(.A(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n211_), .C1(new_n212_), .C2(KEYINPUT3), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n214_), .B(KEYINPUT79), .C1(G141gat), .C2(G148gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT2), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n216_), .A2(KEYINPUT80), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT80), .B1(new_n216_), .B2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n209_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n217_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n208_), .B1(new_n207_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT1), .B1(new_n205_), .B2(new_n206_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n227_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n204_), .B1(new_n224_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G197gat), .B(G204gat), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT21), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G197gat), .B(G204gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT21), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT83), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G218gat), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n242_), .A2(G211gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(G211gat), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n243_), .A2(new_n244_), .A3(KEYINPUT83), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n235_), .B(new_n238_), .C1(new_n241_), .C2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT83), .B1(new_n243_), .B2(new_n244_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n239_), .A2(new_n240_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT21), .A4(new_n234_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n203_), .B1(new_n233_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n216_), .A2(new_n221_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n216_), .A2(KEYINPUT80), .A3(new_n221_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n231_), .B1(new_n257_), .B2(new_n209_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n202_), .B(new_n252_), .C1(new_n258_), .C2(new_n204_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n251_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G78gat), .B(G106gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n251_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n258_), .B2(new_n204_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n224_), .A2(new_n204_), .A3(new_n232_), .A4(new_n267_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G22gat), .B(G50gat), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n268_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n224_), .A2(new_n232_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n266_), .B1(new_n274_), .B2(KEYINPUT29), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n271_), .B1(new_n275_), .B2(new_n269_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT86), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n265_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n265_), .B2(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT85), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n272_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n275_), .A2(new_n271_), .A3(new_n269_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(KEYINPUT82), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT84), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n262_), .A2(new_n289_), .A3(new_n264_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n251_), .A2(new_n259_), .A3(KEYINPUT84), .A4(new_n263_), .ZN(new_n291_));
  AND4_X1   g090(.A1(new_n282_), .A2(new_n288_), .A3(new_n290_), .A4(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n291_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n282_), .B1(new_n294_), .B2(new_n290_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n281_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT25), .B(G183gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT26), .B(G190gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G169gat), .ZN(new_n300_));
  INV_X1    g099(.A(G176gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT75), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(G169gat), .B2(G176gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n302_), .A2(new_n304_), .A3(KEYINPUT24), .A4(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT76), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n299_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT24), .B1(new_n302_), .B2(new_n304_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n308_), .A2(new_n310_), .A3(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n312_), .B(KEYINPUT23), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(G183gat), .B2(G190gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n300_), .A2(new_n301_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT22), .B(G169gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n320_), .B2(new_n301_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT30), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT77), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n323_), .B(KEYINPUT30), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G71gat), .B(G99gat), .ZN(new_n330_));
  INV_X1    g129(.A(G43gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G227gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(G15gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n332_), .B(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(new_n329_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n339_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n340_), .A2(KEYINPUT78), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT78), .B1(new_n340_), .B2(new_n341_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT31), .ZN(new_n345_));
  OR3_X1    g144(.A1(new_n327_), .A2(new_n328_), .A3(new_n336_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n337_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n337_), .B2(new_n346_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n296_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n337_), .A2(new_n346_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n345_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n337_), .A2(new_n346_), .A3(new_n345_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n355_), .B(new_n281_), .C1(new_n292_), .C2(new_n295_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n250_), .B1(new_n322_), .B2(new_n316_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT19), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT20), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OR3_X1    g161(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n306_), .A2(new_n317_), .A3(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT26), .B(G190gat), .Z(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT87), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT87), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n298_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n297_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n322_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n362_), .B1(new_n371_), .B2(new_n252_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT88), .B1(new_n358_), .B2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n323_), .A2(new_n252_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n364_), .A2(new_n369_), .B1(new_n321_), .B2(new_n318_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT20), .B1(new_n250_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n360_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n323_), .A2(new_n252_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n250_), .A2(new_n375_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .A4(new_n362_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n373_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G8gat), .B(G36gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n382_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n382_), .A2(new_n388_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT27), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n371_), .B2(new_n252_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n360_), .B1(new_n358_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT97), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT97), .B(new_n360_), .C1(new_n358_), .C2(new_n396_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n374_), .A2(new_n376_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n399_), .B(new_n400_), .C1(new_n360_), .C2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n388_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(KEYINPUT27), .A3(new_n389_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n393_), .A2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G1gat), .B(G29gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G57gat), .B(G85gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT91), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n209_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n415_));
  OAI22_X1  g214(.A1(new_n415_), .A2(new_n231_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT92), .B(KEYINPUT4), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n340_), .A2(new_n341_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n224_), .A2(new_n419_), .A3(new_n232_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(KEYINPUT4), .C1(new_n258_), .C2(new_n344_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n416_), .A2(KEYINPUT90), .A3(KEYINPUT4), .A4(new_n420_), .ZN(new_n424_));
  AOI211_X1 g223(.A(new_n413_), .B(new_n418_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n416_), .A2(new_n420_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(G225gat), .B2(G233gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n410_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n418_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n412_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n427_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n410_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n405_), .A2(new_n434_), .ZN(new_n435_));
  AOI211_X1 g234(.A(new_n427_), .B(new_n410_), .C1(new_n429_), .C2(new_n412_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT33), .B1(new_n436_), .B2(KEYINPUT94), .ZN(new_n437_));
  INV_X1    g236(.A(new_n391_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT94), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n433_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n426_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n432_), .B1(new_n442_), .B2(new_n412_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n429_), .A2(KEYINPUT95), .A3(new_n411_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT95), .B1(new_n429_), .B2(new_n411_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n437_), .A2(new_n438_), .A3(new_n441_), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n387_), .A2(KEYINPUT32), .ZN(new_n448_));
  AND4_X1   g247(.A1(new_n381_), .A2(new_n373_), .A3(new_n377_), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n402_), .B2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n432_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n436_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT98), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n434_), .A2(KEYINPUT98), .A3(new_n451_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n447_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n349_), .B(new_n281_), .C1(new_n292_), .C2(new_n295_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n357_), .A2(new_n435_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G85gat), .B(G92gat), .Z(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT10), .B(G99gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT64), .B(G106gat), .ZN(new_n463_));
  AOI22_X1  g262(.A1(KEYINPUT9), .A2(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT9), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G85gat), .A3(G92gat), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT65), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G29gat), .B(G36gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT67), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT7), .ZN(new_n479_));
  NOR3_X1   g278(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n466_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n480_), .A2(new_n479_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n478_), .B(new_n461_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n461_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n472_), .A2(new_n475_), .A3(new_n483_), .A4(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n470_), .A2(new_n471_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT65), .B1(new_n464_), .B2(new_n469_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n485_), .B(new_n483_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n475_), .B(KEYINPUT15), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G232gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT34), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT35), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(KEYINPUT35), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT70), .Z(new_n498_));
  AND4_X1   g297(.A1(new_n486_), .A2(new_n491_), .A3(new_n496_), .A4(new_n498_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n489_), .A2(new_n490_), .B1(new_n495_), .B2(new_n494_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n500_), .B2(new_n486_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT71), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G190gat), .B(G218gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(G134gat), .B(G162gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n506_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n502_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  OAI221_X1 g310(.A(KEYINPUT71), .B1(new_n511_), .B2(new_n507_), .C1(new_n499_), .C2(new_n501_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n460_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515_));
  INV_X1    g314(.A(G1gat), .ZN(new_n516_));
  INV_X1    g315(.A(G8gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT14), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G1gat), .B(G8gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(new_n475_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n521_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n490_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n475_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n524_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  OAI22_X1  g327(.A1(new_n523_), .A2(new_n524_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT74), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n529_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G127gat), .B(G155gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT16), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G183gat), .B(G211gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n543_));
  XOR2_X1   g342(.A(G71gat), .B(G78gat), .Z(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n543_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n521_), .B(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n540_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT17), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n550_), .B2(new_n540_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n547_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n489_), .A2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n472_), .A2(new_n483_), .A3(new_n485_), .A4(new_n547_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(KEYINPUT12), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n489_), .A2(new_n561_), .A3(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n558_), .A2(new_n559_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(G230gat), .A3(G233gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G120gat), .B(G148gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n568_), .A2(new_n570_), .A3(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(KEYINPUT13), .A3(new_n579_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n514_), .A2(new_n536_), .A3(new_n556_), .A4(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n434_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G1gat), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT101), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT38), .ZN(new_n589_));
  INV_X1    g388(.A(new_n356_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n287_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT82), .B1(new_n285_), .B2(new_n286_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n290_), .B(new_n291_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT85), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n294_), .A2(new_n282_), .A3(new_n290_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n355_), .B1(new_n596_), .B2(new_n281_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n435_), .B1(new_n590_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n457_), .A2(new_n459_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n536_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT99), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n582_), .A2(new_n583_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(KEYINPUT72), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(KEYINPUT72), .ZN(new_n606_));
  AOI211_X1 g405(.A(new_n605_), .B(new_n606_), .C1(new_n510_), .C2(new_n512_), .ZN(new_n607_));
  AND4_X1   g406(.A1(KEYINPUT72), .A2(new_n510_), .A3(new_n604_), .A4(new_n512_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n556_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n603_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n602_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n586_), .A2(G1gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(KEYINPUT100), .A3(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n602_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n619_), .B2(new_n589_), .ZN(new_n621_));
  AOI211_X1 g420(.A(KEYINPUT102), .B(KEYINPUT38), .C1(new_n615_), .C2(new_n618_), .ZN(new_n622_));
  OAI221_X1 g421(.A(new_n588_), .B1(new_n589_), .B2(new_n619_), .C1(new_n621_), .C2(new_n622_), .ZN(G1324gat));
  INV_X1    g422(.A(new_n405_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G8gat), .B1(new_n585_), .B2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT39), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n613_), .A2(new_n517_), .A3(new_n405_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g428(.A(G15gat), .B1(new_n585_), .B2(new_n349_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT41), .Z(new_n631_));
  NAND3_X1  g430(.A1(new_n613_), .A2(new_n334_), .A3(new_n355_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(new_n296_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G22gat), .B1(new_n585_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT42), .ZN(new_n636_));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n613_), .A2(new_n637_), .A3(new_n296_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT103), .Z(G1327gat));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n600_), .B2(new_n610_), .ZN(new_n642_));
  AOI211_X1 g441(.A(KEYINPUT43), .B(new_n609_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n584_), .A2(new_n536_), .A3(new_n611_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(KEYINPUT104), .A3(new_n647_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(KEYINPUT104), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(KEYINPUT104), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n649_), .B(new_n650_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n586_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n513_), .A2(new_n611_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT105), .Z(new_n655_));
  AND2_X1   g454(.A1(new_n584_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n602_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n586_), .A2(G29gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT106), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n653_), .B1(new_n658_), .B2(new_n660_), .ZN(G1328gat));
  NOR2_X1   g460(.A1(new_n624_), .A2(G36gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n602_), .A2(new_n656_), .A3(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT45), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n624_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G36gat), .B1(new_n665_), .B2(KEYINPUT107), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n667_), .B(new_n624_), .C1(new_n648_), .C2(new_n651_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  OAI221_X1 g471(.A(new_n664_), .B1(new_n670_), .B2(KEYINPUT46), .C1(new_n666_), .C2(new_n668_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1329gat));
  OAI21_X1  g473(.A(G43gat), .B1(new_n652_), .B2(new_n349_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n657_), .A2(new_n331_), .A3(new_n355_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1330gat));
  OR3_X1    g478(.A1(new_n658_), .A2(G50gat), .A3(new_n634_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT109), .B1(new_n652_), .B2(new_n634_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G50gat), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n652_), .A2(KEYINPUT109), .A3(new_n634_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1331gat));
  NAND4_X1  g483(.A1(new_n514_), .A2(new_n535_), .A3(new_n556_), .A4(new_n603_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G57gat), .B1(new_n685_), .B2(new_n586_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n584_), .A2(new_n460_), .A3(new_n536_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n609_), .A3(new_n556_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n586_), .A2(G57gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(G1332gat));
  OAI21_X1  g489(.A(G64gat), .B1(new_n685_), .B2(new_n624_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT48), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n624_), .A2(G64gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n688_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT110), .ZN(G1333gat));
  OAI21_X1  g494(.A(G71gat), .B1(new_n685_), .B2(new_n349_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT49), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n349_), .A2(G71gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n688_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT111), .Z(G1334gat));
  OAI21_X1  g499(.A(G78gat), .B1(new_n685_), .B2(new_n634_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT50), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n634_), .A2(G78gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n688_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT112), .ZN(G1335gat));
  INV_X1    g504(.A(G85gat), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT113), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n687_), .A2(new_n707_), .A3(new_n655_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n687_), .B2(new_n655_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n710_), .B2(new_n586_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT114), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n712_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n460_), .B2(new_n609_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n600_), .A2(new_n641_), .A3(new_n610_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI211_X1 g516(.A(new_n536_), .B(new_n556_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n586_), .A2(new_n706_), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n713_), .A2(new_n714_), .B1(new_n719_), .B2(new_n720_), .ZN(G1336gat));
  AND2_X1   g520(.A1(new_n719_), .A2(new_n405_), .ZN(new_n722_));
  INV_X1    g521(.A(G92gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n405_), .A2(new_n723_), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n722_), .A2(new_n723_), .B1(new_n710_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT115), .ZN(G1337gat));
  AND2_X1   g525(.A1(new_n719_), .A2(new_n355_), .ZN(new_n727_));
  INV_X1    g526(.A(G99gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n355_), .A2(new_n462_), .ZN(new_n729_));
  OAI22_X1  g528(.A1(new_n727_), .A2(new_n728_), .B1(new_n710_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g530(.A(new_n296_), .B(new_n718_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT117), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT117), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n717_), .A2(new_n735_), .A3(new_n296_), .A4(new_n718_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n733_), .A2(G106gat), .A3(new_n734_), .A4(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT119), .ZN(new_n738_));
  INV_X1    g537(.A(G106gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n732_), .B2(KEYINPUT117), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT119), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n734_), .A4(new_n736_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n736_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n734_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT120), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT120), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n747_), .B(new_n734_), .C1(new_n740_), .C2(new_n736_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n743_), .A2(new_n746_), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n710_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n296_), .A2(new_n463_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n750_), .A2(KEYINPUT116), .A3(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT53), .B1(new_n749_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n744_), .A2(new_n745_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n747_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n744_), .A2(KEYINPUT120), .A3(new_n745_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n759_), .A2(new_n738_), .A3(new_n742_), .A4(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n754_), .A4(new_n755_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n757_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n612_), .A2(new_n765_), .A3(new_n535_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n612_), .B2(new_n535_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n513_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n579_), .A2(new_n536_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n563_), .A2(new_n565_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT68), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n563_), .A2(new_n565_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n563_), .A2(new_n565_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(KEYINPUT55), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n577_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n770_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n529_), .A2(new_n533_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n524_), .B(new_n526_), .C1(new_n521_), .C2(new_n475_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n534_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(KEYINPUT121), .B2(new_n788_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n788_), .A2(KEYINPUT121), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n580_), .A2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n769_), .B1(new_n784_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT122), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT57), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n782_), .A2(new_n783_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n579_), .A2(new_n536_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n580_), .A2(new_n791_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(KEYINPUT122), .A3(new_n769_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n795_), .A2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n800_), .A2(KEYINPUT124), .A3(KEYINPUT57), .A4(new_n769_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n579_), .A2(new_n791_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT123), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT123), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n579_), .A2(new_n806_), .A3(new_n791_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n805_), .A2(new_n807_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n609_), .B1(new_n808_), .B2(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n805_), .A2(new_n807_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n796_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n809_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT57), .B(new_n769_), .C1(new_n784_), .C2(new_n792_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n802_), .A2(new_n803_), .A3(new_n814_), .A4(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n768_), .B1(new_n818_), .B2(new_n611_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n405_), .A2(new_n586_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n356_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n819_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n825_), .A2(G113gat), .A3(new_n535_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n823_), .A2(KEYINPUT59), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT125), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n795_), .A2(new_n801_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n814_), .A2(new_n803_), .A3(new_n817_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n828_), .B(new_n611_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n768_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n828_), .B1(new_n818_), .B2(new_n611_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n827_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT59), .B1(new_n819_), .B2(new_n823_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n536_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G113gat), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n826_), .A2(new_n838_), .ZN(G1340gat));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n584_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n824_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n835_), .A2(new_n603_), .A3(new_n836_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n840_), .ZN(G1341gat));
  OR3_X1    g643(.A1(new_n825_), .A2(G127gat), .A3(new_n611_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n835_), .A2(new_n556_), .A3(new_n836_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G127gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1342gat));
  OR3_X1    g647(.A1(new_n825_), .A2(G134gat), .A3(new_n769_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n835_), .A2(new_n610_), .A3(new_n836_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(G134gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1343gat));
  NOR2_X1   g651(.A1(new_n819_), .A2(new_n350_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n536_), .A3(new_n820_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n603_), .A3(new_n820_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g656(.A1(new_n853_), .A2(new_n556_), .A3(new_n820_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  AND4_X1   g659(.A1(G162gat), .A2(new_n853_), .A3(new_n610_), .A4(new_n820_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n611_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n832_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n863_), .A2(new_n597_), .A3(new_n513_), .A4(new_n820_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n206_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT126), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(KEYINPUT126), .A3(new_n206_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n861_), .B1(new_n867_), .B2(new_n868_), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n624_), .A2(new_n434_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n355_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n296_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n536_), .B(new_n872_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G169gat), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n862_), .A2(KEYINPUT125), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n832_), .A3(new_n831_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n879_), .A2(new_n536_), .A3(new_n320_), .A4(new_n872_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n877_), .A3(new_n880_), .ZN(G1348gat));
  NAND2_X1  g680(.A1(new_n863_), .A2(new_n634_), .ZN(new_n882_));
  NOR4_X1   g681(.A1(new_n882_), .A2(new_n301_), .A3(new_n584_), .A4(new_n871_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n879_), .A2(new_n603_), .A3(new_n872_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n301_), .B2(new_n884_), .ZN(G1349gat));
  NOR2_X1   g684(.A1(new_n611_), .A2(new_n297_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n872_), .B(new_n886_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(G183gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n870_), .A2(new_n355_), .A3(new_n556_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n882_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n887_), .A2(new_n888_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1350gat));
  NAND2_X1  g694(.A1(new_n879_), .A2(new_n872_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G190gat), .B1(new_n896_), .B2(new_n609_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n513_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n896_), .B2(new_n898_), .ZN(G1351gat));
  NAND3_X1  g698(.A1(new_n853_), .A2(new_n536_), .A3(new_n870_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g700(.A1(new_n853_), .A2(new_n603_), .A3(new_n870_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  AND3_X1   g702(.A1(new_n853_), .A2(new_n556_), .A3(new_n870_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT63), .B(G211gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n904_), .B2(new_n907_), .ZN(G1354gat));
  NAND4_X1  g707(.A1(new_n853_), .A2(new_n242_), .A3(new_n513_), .A4(new_n870_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n853_), .A2(new_n610_), .A3(new_n870_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n242_), .ZN(G1355gat));
endmodule


