//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR3_X1   g010(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT66), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT65), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  AND3_X1   g018(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n210_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n213_), .A2(new_n218_), .A3(new_n222_), .A4(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G85gat), .B(G92gat), .Z(new_n230_));
  AND2_X1   g029(.A1(new_n230_), .A2(KEYINPUT8), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(KEYINPUT10), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT10), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G99gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(G106gat), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n216_), .A2(new_n217_), .ZN(new_n236_));
  INV_X1    g035(.A(G85gat), .ZN(new_n237_));
  INV_X1    g036(.A(G92gat), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT9), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n235_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n230_), .A2(KEYINPUT9), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n229_), .A2(new_n231_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n226_), .A2(new_n216_), .A3(new_n217_), .A4(new_n210_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n220_), .A2(new_n221_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n246_), .A2(KEYINPUT64), .A3(new_n210_), .A4(new_n226_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n247_), .A3(new_n230_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT8), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n209_), .B1(new_n242_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n202_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT12), .B1(new_n251_), .B2(new_n202_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G230gat), .ZN(new_n256_));
  INV_X1    g055(.A(G233gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n242_), .A2(new_n250_), .A3(new_n209_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n202_), .B(KEYINPUT12), .C1(new_n251_), .C2(new_n252_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n255_), .A2(new_n259_), .A3(new_n260_), .A4(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n260_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n258_), .B1(new_n263_), .B2(new_n251_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G176gat), .B(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n262_), .A2(new_n264_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n270_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT13), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT71), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n262_), .A2(new_n264_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n269_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n271_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(KEYINPUT13), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT70), .B1(new_n278_), .B2(KEYINPUT13), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT13), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n277_), .A2(new_n283_), .A3(new_n284_), .A4(new_n271_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G190gat), .B(G218gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(G134gat), .B(G162gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT36), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT36), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n242_), .A2(new_n250_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G29gat), .B(G36gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G43gat), .B(G50gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n293_), .B1(new_n294_), .B2(new_n298_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n242_), .A2(new_n250_), .A3(KEYINPUT73), .A4(new_n297_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT34), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT35), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n297_), .B(KEYINPUT15), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n294_), .A2(new_n307_), .A3(KEYINPUT72), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT72), .B1(new_n294_), .B2(new_n307_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n301_), .B(new_n306_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n304_), .A2(new_n305_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n310_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n308_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n312_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n306_), .A4(new_n301_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n292_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n291_), .B1(new_n318_), .B2(new_n290_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n317_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT74), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n321_), .B(new_n291_), .C1(new_n318_), .C2(new_n290_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(KEYINPUT75), .A2(KEYINPUT37), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT76), .B(G22gat), .ZN(new_n328_));
  INV_X1    g127(.A(G15gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G1gat), .ZN(new_n331_));
  INV_X1    g130(.A(G8gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT14), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G1gat), .B(G8gat), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(new_n209_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G231gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT17), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G183gat), .B(G211gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G127gat), .B(G155gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n341_), .A2(new_n342_), .A3(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(KEYINPUT17), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n341_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT75), .B(KEYINPUT37), .Z(new_n353_));
  NAND3_X1  g152(.A1(new_n323_), .A2(new_n324_), .A3(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n287_), .A2(new_n327_), .A3(new_n352_), .A4(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(KEYINPUT78), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n338_), .A2(new_n298_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n297_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n359_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(G229gat), .A4(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n358_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n338_), .A2(new_n307_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G229gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT80), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G141gat), .ZN(new_n369_));
  INV_X1    g168(.A(G197gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT81), .B(G169gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  NAND3_X1  g172(.A1(new_n363_), .A2(new_n368_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n357_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(KEYINPUT82), .A3(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT19), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT94), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT21), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G211gat), .B(G218gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n384_), .B2(new_n383_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT95), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(KEYINPUT95), .A3(new_n389_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT93), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n383_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(new_n386_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n388_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G183gat), .A2(G190gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT23), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT85), .B(KEYINPUT23), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n403_), .B2(new_n400_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n401_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n400_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(new_n402_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT88), .B1(new_n411_), .B2(new_n406_), .ZN(new_n412_));
  INV_X1    g211(.A(G176gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(KEYINPUT22), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G169gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT22), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(G169gat), .B2(G176gat), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n419_), .B(new_n414_), .C1(G169gat), .C2(new_n418_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n408_), .A2(new_n412_), .A3(new_n416_), .A4(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(G169gat), .B2(G176gat), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n423_), .A2(KEYINPUT84), .ZN(new_n424_));
  NOR3_X1   g223(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n423_), .B2(KEYINPUT84), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT23), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n410_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n402_), .B2(new_n410_), .ZN(new_n429_));
  INV_X1    g228(.A(G190gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT83), .B1(new_n430_), .B2(KEYINPUT26), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT25), .B(G183gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT26), .B(G190gat), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n431_), .B(new_n432_), .C1(new_n433_), .C2(KEYINPUT83), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n424_), .A2(new_n426_), .A3(new_n429_), .A4(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n421_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n399_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n411_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n433_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n432_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n429_), .A2(new_n407_), .B1(G169gat), .B2(G176gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT22), .B(G169gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n413_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n392_), .A2(new_n393_), .B1(new_n388_), .B2(new_n397_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n438_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n437_), .B1(new_n449_), .B2(KEYINPUT99), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT99), .ZN(new_n451_));
  AOI211_X1 g250(.A(new_n451_), .B(new_n438_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n382_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT97), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n442_), .A2(new_n446_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n399_), .A2(KEYINPUT97), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n438_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n382_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n448_), .A2(new_n435_), .A3(new_n421_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n453_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G8gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(G92gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT18), .B(G64gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n462_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n449_), .A2(new_n459_), .A3(new_n437_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n458_), .A2(new_n460_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n466_), .B(new_n469_), .C1(new_n470_), .C2(new_n459_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n459_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n469_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n467_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n472_), .A2(KEYINPUT27), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G225gat), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G155gat), .A2(G162gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n481_), .B1(new_n482_), .B2(KEYINPUT1), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(KEYINPUT1), .ZN(new_n484_));
  OR2_X1    g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT1), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n486_), .A2(KEYINPUT90), .A3(G155gat), .A4(G162gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .A4(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(G141gat), .A2(G148gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G141gat), .A2(G148gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT91), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G141gat), .A2(G148gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT2), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n490_), .B(new_n496_), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n495_), .A2(new_n497_), .A3(KEYINPUT92), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT92), .B1(new_n495_), .B2(new_n497_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n482_), .A4(new_n485_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G127gat), .B(G134gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G113gat), .B(G120gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n506_), .A2(KEYINPUT4), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n492_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(KEYINPUT4), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n480_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n506_), .A2(new_n508_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n480_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G57gat), .B(G85gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G1gat), .B(G29gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n514_), .A2(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n510_), .A2(new_n513_), .A3(new_n519_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G78gat), .B(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n501_), .A2(KEYINPUT29), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G228gat), .A2(G233gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n399_), .A3(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n528_));
  AOI21_X1  g327(.A(new_n448_), .B1(new_n501_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n530_), .A2(G22gat), .ZN(new_n531_));
  INV_X1    g330(.A(G22gat), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n527_), .B(new_n532_), .C1(new_n526_), .C2(new_n529_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n524_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n501_), .A2(KEYINPUT29), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(KEYINPUT28), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(KEYINPUT28), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G50gat), .ZN(new_n540_));
  INV_X1    g339(.A(G50gat), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n541_), .A3(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n530_), .A2(G22gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n524_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n533_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n535_), .A2(new_n540_), .A3(new_n542_), .A4(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n542_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n533_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n544_), .B1(new_n543_), .B2(new_n533_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G15gat), .B(G43gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G227gat), .A2(G233gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n421_), .A2(new_n555_), .A3(new_n435_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n555_), .B1(new_n421_), .B2(new_n435_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n505_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n504_), .A3(new_n556_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n554_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G71gat), .B(G99gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(new_n561_), .A3(new_n554_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n566_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n567_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n570_), .B2(new_n562_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n546_), .A2(new_n550_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n479_), .B(new_n523_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n572_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT100), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n466_), .A2(KEYINPUT32), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n462_), .B2(new_n580_), .ZN(new_n581_));
  AOI211_X1 g380(.A(KEYINPUT100), .B(new_n579_), .C1(new_n453_), .C2(new_n461_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n473_), .A2(new_n474_), .A3(new_n580_), .ZN(new_n583_));
  NOR4_X1   g382(.A1(new_n523_), .A2(new_n581_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n512_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n511_), .A2(new_n480_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n519_), .B1(new_n587_), .B2(KEYINPUT33), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT33), .B(new_n519_), .C1(new_n510_), .C2(new_n513_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n510_), .A2(new_n513_), .A3(KEYINPUT33), .ZN(new_n591_));
  NOR4_X1   g390(.A1(new_n476_), .A2(new_n588_), .A3(new_n590_), .A4(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n577_), .B1(new_n584_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n575_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n355_), .A2(KEYINPUT78), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n356_), .A2(new_n380_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT102), .Z(new_n597_));
  INV_X1    g396(.A(new_n523_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n331_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n594_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n325_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n351_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n380_), .A3(new_n287_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G1gat), .B1(new_n605_), .B2(new_n523_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n599_), .A2(new_n600_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n601_), .A2(new_n606_), .A3(new_n607_), .ZN(G1324gat));
  OAI21_X1  g407(.A(G8gat), .B1(new_n605_), .B2(new_n479_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT39), .ZN(new_n610_));
  INV_X1    g409(.A(new_n479_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n597_), .A2(new_n332_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n610_), .A2(KEYINPUT40), .A3(new_n612_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1325gat));
  OAI21_X1  g416(.A(G15gat), .B1(new_n605_), .B2(new_n572_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT41), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n597_), .A2(new_n329_), .A3(new_n576_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1326gat));
  NAND2_X1  g420(.A1(new_n546_), .A2(new_n550_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G22gat), .B1(new_n605_), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT42), .ZN(new_n624_));
  INV_X1    g423(.A(new_n622_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n597_), .A2(new_n532_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(G1327gat));
  NAND2_X1  g426(.A1(new_n287_), .A2(new_n380_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(new_n352_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n594_), .A3(new_n603_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT103), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n629_), .A2(new_n594_), .A3(new_n632_), .A4(new_n603_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n598_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n327_), .A2(new_n354_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n594_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n594_), .B2(new_n637_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n629_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT44), .B(new_n629_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n598_), .A2(G29gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n635_), .B1(new_n644_), .B2(new_n645_), .ZN(G1328gat));
  NAND3_X1  g445(.A1(new_n642_), .A2(new_n611_), .A3(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G36gat), .ZN(new_n648_));
  INV_X1    g447(.A(G36gat), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n631_), .A2(new_n649_), .A3(new_n611_), .A4(new_n633_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT104), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT45), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(KEYINPUT104), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n648_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI221_X1 g457(.A(new_n648_), .B1(KEYINPUT105), .B2(KEYINPUT46), .C1(new_n654_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1329gat));
  AND2_X1   g459(.A1(new_n634_), .A2(new_n576_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(G43gat), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n642_), .A2(G43gat), .A3(new_n576_), .A4(new_n643_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(KEYINPUT106), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(KEYINPUT106), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT47), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n668_), .B(new_n662_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1330gat));
  NAND3_X1  g469(.A1(new_n634_), .A2(new_n541_), .A3(new_n625_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n642_), .A2(new_n625_), .A3(new_n643_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT107), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n642_), .A2(new_n674_), .A3(new_n625_), .A4(new_n643_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(G50gat), .A3(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT108), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT108), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n671_), .B1(new_n677_), .B2(new_n678_), .ZN(G1331gat));
  INV_X1    g478(.A(new_n380_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n287_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n604_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT110), .B1(new_n523_), .B2(new_n683_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n682_), .A2(KEYINPUT110), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n684_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n323_), .A2(new_n324_), .A3(new_n353_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n326_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n687_), .A2(new_n689_), .A3(new_n351_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n681_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT109), .Z(new_n692_));
  NOR2_X1   g491(.A1(new_n602_), .A2(new_n380_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n695_), .A3(new_n598_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n685_), .B1(new_n696_), .B2(new_n683_), .ZN(G1332gat));
  INV_X1    g496(.A(G64gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n682_), .B2(new_n611_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT48), .Z(new_n700_));
  NAND2_X1  g499(.A1(new_n611_), .A2(new_n698_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n694_), .B2(new_n701_), .ZN(G1333gat));
  INV_X1    g501(.A(G71gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n682_), .B2(new_n576_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT49), .Z(new_n705_));
  NAND3_X1  g504(.A1(new_n695_), .A2(new_n703_), .A3(new_n576_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1334gat));
  INV_X1    g506(.A(G78gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n682_), .B2(new_n625_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT50), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n695_), .A2(new_n708_), .A3(new_n625_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1335gat));
  NOR3_X1   g511(.A1(new_n287_), .A2(new_n380_), .A3(new_n352_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n594_), .A2(new_n603_), .A3(new_n713_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n714_), .A2(G85gat), .A3(new_n523_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n598_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n715_), .B1(new_n718_), .B2(G85gat), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT111), .Z(G1336gat));
  INV_X1    g519(.A(new_n714_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G92gat), .B1(new_n721_), .B2(new_n611_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n611_), .A2(G92gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT112), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n717_), .B2(new_n724_), .ZN(G1337gat));
  OAI21_X1  g524(.A(G99gat), .B1(new_n716_), .B2(new_n572_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n572_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n721_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n726_), .B(new_n728_), .C1(KEYINPUT113), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(KEYINPUT51), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n730_), .B(new_n732_), .Z(G1338gat));
  OAI21_X1  g532(.A(G106gat), .B1(new_n716_), .B2(new_n622_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT52), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n721_), .A2(new_n225_), .A3(new_n625_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1339gat));
  OAI21_X1  g538(.A(KEYINPUT115), .B1(new_n355_), .B2(new_n380_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n690_), .A2(new_n741_), .A3(new_n680_), .A4(new_n287_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT54), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n742_), .A3(KEYINPUT54), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n255_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n258_), .A2(KEYINPUT116), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT55), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n749_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n253_), .A2(new_n254_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n261_), .A2(new_n260_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT55), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n751_), .B1(new_n756_), .B2(new_n262_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT117), .B1(new_n757_), .B2(new_n270_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n748_), .B2(new_n752_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n262_), .ZN(new_n762_));
  OAI22_X1  g561(.A1(new_n761_), .A2(new_n762_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n269_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n758_), .A2(new_n759_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT118), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(KEYINPUT56), .A3(new_n269_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n758_), .A2(new_n769_), .A3(new_n759_), .A4(new_n765_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n768_), .A3(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n680_), .A2(new_n272_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n361_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n373_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n364_), .A2(new_n365_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT119), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT119), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n364_), .A2(new_n778_), .A3(new_n365_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n774_), .B(new_n775_), .C1(new_n780_), .C2(new_n367_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n374_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n278_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT120), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n785_), .A3(new_n278_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n773_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT57), .A3(new_n325_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n763_), .A2(new_n269_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n759_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT121), .A3(new_n768_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n794_), .A3(new_n759_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n793_), .A2(new_n271_), .A3(new_n782_), .A4(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n797_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n637_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n787_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n603_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n790_), .A2(new_n800_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n747_), .B1(new_n351_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n574_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n611_), .A2(new_n523_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n805_), .A2(new_n806_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n380_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n804_), .A2(new_n351_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n745_), .A2(new_n746_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(new_n574_), .A3(new_n807_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n813_), .A2(KEYINPUT59), .A3(new_n574_), .A4(new_n807_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n680_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n810_), .B1(new_n818_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g618(.A(G120gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n287_), .B2(KEYINPUT60), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n809_), .B(new_n821_), .C1(KEYINPUT60), .C2(new_n820_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n287_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n820_), .ZN(G1341gat));
  AOI21_X1  g623(.A(G127gat), .B1(new_n809_), .B2(new_n352_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n816_), .A2(new_n817_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n352_), .A2(G127gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT122), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n825_), .B1(new_n826_), .B2(new_n828_), .ZN(G1342gat));
  AOI21_X1  g628(.A(G134gat), .B1(new_n809_), .B2(new_n603_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n637_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n832_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g632(.A(new_n573_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n805_), .A2(new_n834_), .A3(new_n808_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n380_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n681_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g638(.A1(new_n835_), .A2(new_n352_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT61), .B(G155gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT123), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n840_), .B(new_n843_), .ZN(G1346gat));
  AOI21_X1  g643(.A(G162gat), .B1(new_n835_), .B2(new_n603_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n637_), .A2(G162gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n835_), .B2(new_n846_), .ZN(G1347gat));
  NOR2_X1   g646(.A1(new_n479_), .A2(new_n598_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n813_), .A2(new_n380_), .A3(new_n574_), .A4(new_n848_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n850_));
  AND3_X1   g649(.A1(new_n849_), .A2(G169gat), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n849_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n852_), .B2(new_n444_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(G169gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n851_), .B1(new_n853_), .B2(new_n854_), .ZN(G1348gat));
  NAND3_X1  g654(.A1(new_n813_), .A2(new_n574_), .A3(new_n848_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n856_), .A2(new_n287_), .B1(KEYINPUT125), .B2(new_n413_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n848_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n805_), .A2(new_n806_), .A3(new_n858_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT125), .B(G176gat), .Z(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n681_), .A3(new_n860_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n857_), .A2(new_n861_), .ZN(G1349gat));
  INV_X1    g661(.A(KEYINPUT126), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n859_), .A2(new_n863_), .A3(new_n441_), .A4(new_n352_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n813_), .A2(new_n574_), .A3(new_n352_), .A4(new_n848_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT126), .B1(new_n865_), .B2(new_n432_), .ZN(new_n866_));
  INV_X1    g665(.A(G183gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n864_), .A2(new_n866_), .A3(new_n868_), .ZN(G1350gat));
  NAND3_X1  g668(.A1(new_n859_), .A2(new_n603_), .A3(new_n433_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G190gat), .B1(new_n856_), .B2(new_n831_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1351gat));
  NOR3_X1   g671(.A1(new_n805_), .A2(new_n834_), .A3(new_n858_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n873_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n380_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT127), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n813_), .A2(new_n380_), .A3(new_n573_), .A4(new_n848_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n370_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n370_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n874_), .A2(new_n877_), .A3(new_n878_), .ZN(G1352gat));
  NAND2_X1  g678(.A1(new_n873_), .A2(new_n681_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g680(.A(KEYINPUT63), .B(G211gat), .Z(new_n882_));
  AND3_X1   g681(.A1(new_n873_), .A2(new_n352_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n873_), .A2(new_n352_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1354gat));
  AOI21_X1  g685(.A(G218gat), .B1(new_n873_), .B2(new_n603_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n637_), .A2(G218gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n873_), .B2(new_n888_), .ZN(G1355gat));
endmodule


