//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_;
  XNOR2_X1  g000(.A(KEYINPUT0), .B(G57gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G1gat), .B(G29gat), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT90), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n212_), .A2(new_n213_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n219_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n214_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n218_), .A2(new_n221_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G113gat), .B(G120gat), .Z(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT87), .B(G127gat), .ZN(new_n229_));
  INV_X1    g028(.A(G134gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G127gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n232_), .A2(KEYINPUT87), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(KEYINPUT87), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n233_), .A2(new_n234_), .A3(G134gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n228_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(G134gat), .B1(new_n233_), .B2(new_n234_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n229_), .A2(new_n230_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n227_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n236_), .A2(KEYINPUT88), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT88), .B1(new_n236_), .B2(new_n239_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n226_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n225_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT99), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(KEYINPUT99), .A3(new_n244_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n206_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n242_), .A2(KEYINPUT4), .A3(new_n244_), .ZN(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT98), .B(KEYINPUT4), .Z(new_n251_));
  OAI211_X1 g050(.A(new_n226_), .B(new_n251_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n246_), .A3(new_n252_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n253_), .A2(KEYINPUT100), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(KEYINPUT100), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n249_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G204gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G197gat), .ZN(new_n258_));
  INV_X1    g057(.A(G197gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G204gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(G211gat), .A2(G218gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G211gat), .A2(G218gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n261_), .A2(new_n264_), .A3(KEYINPUT21), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT93), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT93), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n264_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n258_), .A2(new_n260_), .A3(new_n267_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n268_), .A2(new_n264_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n266_), .A2(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G190gat), .ZN(new_n278_));
  INV_X1    g077(.A(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT26), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n278_), .A2(new_n280_), .A3(KEYINPUT96), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT96), .B1(new_n278_), .B2(new_n280_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n276_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(G183gat), .B2(G190gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT23), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n286_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT97), .ZN(new_n292_));
  INV_X1    g091(.A(new_n284_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT24), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(KEYINPUT23), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n287_), .A2(G183gat), .A3(G190gat), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n296_), .A2(new_n297_), .B1(new_n285_), .B2(new_n284_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT97), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n283_), .A2(new_n292_), .A3(new_n295_), .A4(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT22), .B(G169gat), .ZN(new_n302_));
  INV_X1    g101(.A(G176gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n296_), .A2(new_n297_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n304_), .B(new_n294_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n273_), .A2(new_n301_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n261_), .A2(KEYINPUT21), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n309_), .B(new_n271_), .C1(new_n263_), .C2(new_n262_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n270_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n269_), .B1(new_n268_), .B2(new_n264_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n277_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n278_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n298_), .B(new_n295_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT22), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n303_), .B1(new_n319_), .B2(KEYINPUT82), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G169gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n284_), .B1(KEYINPUT82), .B2(new_n319_), .ZN(new_n322_));
  AOI21_X1  g121(.A(G183gat), .B1(new_n314_), .B2(new_n315_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n321_), .B(new_n322_), .C1(new_n305_), .C2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n313_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n308_), .A2(KEYINPUT20), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT19), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n301_), .A2(new_n307_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n313_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n273_), .A2(new_n324_), .A3(new_n318_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n333_), .A2(KEYINPUT20), .A3(new_n329_), .A4(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT18), .B(G64gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G92gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n331_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT33), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n250_), .A2(G225gat), .A3(G233gat), .A4(new_n252_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n242_), .A2(new_n246_), .A3(new_n244_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n344_), .B1(new_n347_), .B2(new_n205_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(KEYINPUT33), .A4(new_n206_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n256_), .A2(new_n343_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n331_), .A2(new_n335_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT32), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(new_n340_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n327_), .A2(new_n329_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n333_), .A2(KEYINPUT20), .A3(new_n330_), .A4(new_n334_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(KEYINPUT32), .A3(new_n339_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n347_), .A2(new_n205_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n206_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n353_), .B(new_n357_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n350_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT30), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n318_), .A2(new_n324_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n318_), .B2(new_n324_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT85), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n325_), .A2(KEYINPUT30), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n318_), .A2(new_n324_), .A3(new_n362_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G15gat), .B(G43gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n372_), .B(new_n375_), .Z(new_n376_));
  NAND3_X1  g175(.A1(new_n365_), .A2(new_n369_), .A3(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n372_), .B(new_n375_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n378_), .B(KEYINPUT85), .C1(new_n364_), .C2(new_n363_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT86), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT31), .ZN(new_n382_));
  INV_X1    g181(.A(new_n241_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n236_), .A2(KEYINPUT88), .A3(new_n239_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT31), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n377_), .A2(new_n388_), .A3(new_n379_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n381_), .A2(KEYINPUT89), .A3(new_n387_), .A4(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n377_), .A2(new_n388_), .A3(new_n379_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n388_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n387_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT89), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n393_), .B2(new_n380_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n390_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n218_), .A2(new_n221_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n224_), .A2(new_n222_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT94), .ZN(new_n403_));
  INV_X1    g202(.A(G228gat), .ZN(new_n404_));
  INV_X1    g203(.A(G233gat), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(KEYINPUT92), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(KEYINPUT92), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  OAI22_X1  g207(.A1(new_n402_), .A2(new_n273_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G78gat), .B(G106gat), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n408_), .B(new_n403_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n313_), .B(new_n412_), .C1(new_n225_), .C2(new_n399_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n409_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n411_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT95), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n409_), .A2(new_n413_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n410_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT95), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n409_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G22gat), .B(G50gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n225_), .B2(new_n399_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n225_), .A2(new_n399_), .A3(new_n425_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n423_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n428_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n430_), .A2(new_n422_), .A3(new_n426_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n416_), .A2(new_n421_), .A3(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n429_), .A2(new_n431_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(new_n419_), .A3(new_n418_), .A4(new_n420_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n361_), .A2(new_n398_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n356_), .A2(new_n340_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n351_), .A2(new_n339_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT27), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT27), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n397_), .A2(new_n443_), .A3(new_n436_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n433_), .A2(new_n435_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT101), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n339_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n342_), .A2(new_n447_), .A3(new_n441_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n331_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT27), .B1(new_n439_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n446_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT101), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n445_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n444_), .B1(new_n453_), .B2(new_n397_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n358_), .A2(new_n359_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n437_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT13), .ZN(new_n457_));
  XOR2_X1   g256(.A(G120gat), .B(G148gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT71), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G176gat), .B(G204gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(KEYINPUT9), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n467_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT9), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT10), .B(G99gat), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n468_), .B(new_n471_), .C1(G106gat), .C2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT7), .ZN(new_n474_));
  INV_X1    g273(.A(G99gat), .ZN(new_n475_));
  INV_X1    g274(.A(G106gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT8), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n473_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n485_));
  AND2_X1   g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n481_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n466_), .A2(new_n467_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n478_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n495_));
  NAND2_X1  g294(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n486_), .A3(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n498_));
  NOR2_X1   g297(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n483_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n497_), .A2(new_n500_), .A3(new_n479_), .A4(new_n477_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n492_), .A2(new_n478_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n494_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G57gat), .ZN(new_n504_));
  INV_X1    g303(.A(G64gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G57gat), .A2(G64gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT11), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G71gat), .B(G78gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT11), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n506_), .A2(new_n512_), .A3(new_n507_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n508_), .A2(new_n510_), .A3(KEYINPUT11), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n491_), .A2(new_n503_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT66), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n491_), .A2(new_n519_), .A3(new_n503_), .A4(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n516_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n501_), .A2(new_n502_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n493_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n489_), .B1(new_n480_), .B2(new_n473_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n522_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT67), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n516_), .B1(new_n491_), .B2(new_n503_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT67), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n521_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G230gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(new_n405_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT68), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n531_), .A2(KEYINPUT68), .A3(new_n533_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n533_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n517_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n529_), .A2(KEYINPUT69), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT69), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT12), .B1(new_n526_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n541_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n463_), .B1(new_n538_), .B2(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n531_), .A2(KEYINPUT68), .A3(new_n533_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT68), .B1(new_n531_), .B2(new_n533_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n546_), .B(new_n463_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n457_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n546_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n463_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(KEYINPUT13), .A3(new_n550_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G8gat), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT76), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G1gat), .A2(G8gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT14), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n560_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G29gat), .B(G36gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G43gat), .ZN(new_n568_));
  INV_X1    g367(.A(G50gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n567_), .A2(G43gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(G43gat), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(G50gat), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT15), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n570_), .A2(KEYINPUT15), .A3(new_n573_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n566_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n566_), .A2(new_n573_), .A3(new_n570_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n579_), .A2(KEYINPUT79), .A3(new_n580_), .A4(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT79), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n560_), .B(new_n564_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n574_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n580_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n583_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n584_), .A2(new_n574_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n578_), .A2(new_n589_), .A3(new_n587_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n582_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G169gat), .B(G197gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT80), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(G113gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(G141gat), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n595_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n582_), .B(new_n597_), .C1(new_n588_), .C2(new_n590_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n557_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n516_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n566_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT17), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n604_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n604_), .A2(new_n612_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n456_), .A2(new_n601_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n576_), .A2(new_n577_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n574_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT34), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(KEYINPUT35), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(KEYINPUT35), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n624_), .A2(KEYINPUT35), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n619_), .A2(new_n626_), .A3(new_n627_), .A4(new_n621_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT72), .B(G190gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(G218gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(G134gat), .B(G162gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT36), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n629_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT74), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n629_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n617_), .B1(new_n635_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n629_), .A2(new_n634_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n617_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n642_), .B(new_n643_), .C1(new_n629_), .C2(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n616_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n455_), .B(KEYINPUT102), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n646_), .A2(G1gat), .A3(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(KEYINPUT38), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT103), .Z(new_n650_));
  NOR2_X1   g449(.A1(new_n635_), .A2(new_n640_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n616_), .A2(new_n652_), .A3(new_n455_), .ZN(new_n653_));
  AOI22_X1  g452(.A1(new_n648_), .A2(KEYINPUT38), .B1(G1gat), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n650_), .A2(new_n654_), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n451_), .A2(new_n452_), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n646_), .A2(G8gat), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n656_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n616_), .A2(new_n652_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n659_), .A2(new_n660_), .A3(G8gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n659_), .B2(G8gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n657_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(KEYINPUT104), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(KEYINPUT104), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(KEYINPUT40), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT40), .B1(new_n664_), .B2(new_n665_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  OR3_X1    g467(.A1(new_n646_), .A2(G15gat), .A3(new_n398_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n616_), .A2(new_n652_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G15gat), .B1(new_n670_), .B2(new_n398_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT105), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(KEYINPUT105), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(KEYINPUT41), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(new_n672_), .B2(new_n673_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n669_), .B1(new_n674_), .B2(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n670_), .B2(new_n436_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n646_), .A2(G22gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n436_), .B2(new_n679_), .ZN(G1327gat));
  AND3_X1   g479(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT101), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT101), .B1(new_n440_), .B2(new_n442_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n397_), .B(new_n436_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n394_), .A2(new_n396_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n448_), .A2(new_n450_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n445_), .A4(new_n390_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n455_), .B1(new_n683_), .B2(new_n686_), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n397_), .B(new_n445_), .C1(new_n350_), .C2(new_n360_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n615_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(new_n651_), .A3(new_n601_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n455_), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n691_), .A2(G29gat), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n615_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  INV_X1    g494(.A(new_n645_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n456_), .B2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n695_), .B(new_n696_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n601_), .B(new_n694_), .C1(new_n697_), .C2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n647_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n689_), .B2(new_n645_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n698_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n705_), .A2(KEYINPUT44), .A3(new_n601_), .A4(new_n694_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n702_), .A2(new_n703_), .A3(new_n706_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n707_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT106), .B1(new_n707_), .B2(G29gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n693_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n691_), .A2(G36gat), .A3(new_n656_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT45), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n702_), .A2(new_n658_), .A3(new_n706_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(G36gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G36gat), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n713_), .B(new_n715_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n711_), .A2(new_n712_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n716_), .A2(G36gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT107), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n716_), .A2(new_n717_), .A3(G36gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n721_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n713_), .A4(new_n715_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n722_), .A2(new_n728_), .ZN(G1329gat));
  NOR3_X1   g528(.A1(new_n691_), .A2(G43gat), .A3(new_n398_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n702_), .A2(new_n397_), .A3(new_n706_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G43gat), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g532(.A1(new_n702_), .A2(new_n445_), .A3(new_n706_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n735_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(G50gat), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n445_), .A2(new_n569_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n691_), .B2(new_n739_), .ZN(G1331gat));
  NAND2_X1  g539(.A1(new_n557_), .A2(new_n600_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n456_), .A2(new_n742_), .A3(new_n615_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n651_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G57gat), .B1(new_n745_), .B2(new_n692_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n743_), .A2(new_n696_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n504_), .A3(new_n703_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT110), .ZN(G1332gat));
  NAND3_X1  g549(.A1(new_n747_), .A2(new_n505_), .A3(new_n658_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n745_), .A2(new_n656_), .ZN(new_n752_));
  OR3_X1    g551(.A1(new_n752_), .A2(KEYINPUT111), .A3(new_n505_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT111), .B1(new_n752_), .B2(new_n505_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(KEYINPUT48), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT48), .B1(new_n753_), .B2(new_n754_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n751_), .B1(new_n755_), .B2(new_n756_), .ZN(G1333gat));
  INV_X1    g556(.A(G71gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n744_), .B2(new_n397_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT49), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n747_), .A2(new_n758_), .A3(new_n397_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1334gat));
  INV_X1    g561(.A(G78gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n744_), .B2(new_n445_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT50), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n747_), .A2(new_n763_), .A3(new_n445_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1335gat));
  NAND3_X1  g566(.A1(new_n705_), .A2(new_n694_), .A3(new_n742_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(KEYINPUT112), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(KEYINPUT112), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(G85gat), .A3(new_n455_), .A4(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n690_), .A2(new_n742_), .A3(new_n651_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n464_), .B1(new_n772_), .B2(new_n647_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1336gat));
  NAND4_X1  g573(.A1(new_n769_), .A2(G92gat), .A3(new_n658_), .A4(new_n770_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n465_), .B1(new_n772_), .B2(new_n656_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1337gat));
  OR3_X1    g576(.A1(new_n772_), .A2(new_n472_), .A3(new_n398_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n769_), .A2(new_n397_), .A3(new_n770_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n475_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT51), .ZN(G1338gat));
  OR2_X1    g580(.A1(new_n768_), .A2(new_n436_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G106gat), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n772_), .A2(G106gat), .A3(new_n436_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT113), .Z(new_n787_));
  NAND3_X1  g586(.A1(new_n782_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g589(.A1(new_n647_), .A2(new_n658_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n397_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT55), .B(new_n541_), .C1(new_n543_), .C2(new_n545_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT117), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n546_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n521_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n533_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n542_), .B1(new_n529_), .B2(KEYINPUT69), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n526_), .A2(new_n544_), .A3(KEYINPUT12), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n540_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(KEYINPUT55), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n795_), .A2(new_n797_), .A3(new_n799_), .A4(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n554_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n554_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n599_), .A2(new_n550_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n599_), .A2(KEYINPUT116), .A3(new_n550_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n806_), .A2(KEYINPUT118), .A3(new_n807_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n811_), .A2(new_n814_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n579_), .A2(new_n587_), .A3(new_n581_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n586_), .A2(new_n580_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n595_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n821_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n822_), .A2(new_n598_), .A3(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n817_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT57), .B1(new_n826_), .B2(new_n652_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n828_), .B(new_n651_), .C1(new_n817_), .C2(new_n825_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n808_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n806_), .A2(KEYINPUT120), .A3(new_n807_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n833_), .A2(new_n810_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n824_), .A2(new_n550_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n831_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n833_), .A2(new_n810_), .A3(new_n834_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(KEYINPUT58), .A3(new_n550_), .A4(new_n824_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n696_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n615_), .B1(new_n830_), .B2(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n555_), .A2(KEYINPUT13), .A3(new_n550_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT13), .B1(new_n555_), .B2(new_n550_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n600_), .A4(new_n615_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n552_), .A2(new_n600_), .A3(new_n556_), .A4(new_n615_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT114), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n848_), .A3(new_n645_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n850_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n846_), .A2(new_n848_), .A3(new_n645_), .A4(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n436_), .B(new_n793_), .C1(new_n841_), .C2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n826_), .A2(new_n652_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n828_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n826_), .A2(KEYINPUT57), .A3(new_n652_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n840_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n694_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n854_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n864_), .A2(KEYINPUT121), .A3(new_n436_), .A4(new_n793_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n857_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G113gat), .B1(new_n866_), .B2(new_n599_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n855_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n445_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT59), .A3(new_n793_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n600_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n867_), .B1(G113gat), .B2(new_n872_), .ZN(G1340gat));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n866_), .B1(KEYINPUT60), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n876_));
  AOI21_X1  g675(.A(G120gat), .B1(new_n557_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n844_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n875_), .A2(new_n877_), .B1(new_n874_), .B2(new_n878_), .ZN(G1341gat));
  AOI211_X1 g678(.A(new_n232_), .B(new_n694_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT121), .B1(new_n870_), .B2(new_n793_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n854_), .B1(new_n861_), .B2(new_n694_), .ZN(new_n882_));
  NOR4_X1   g681(.A1(new_n882_), .A2(new_n856_), .A3(new_n445_), .A4(new_n792_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n615_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n232_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n694_), .B1(new_n857_), .B2(new_n865_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n887_), .B2(G127gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n880_), .B1(new_n886_), .B2(new_n888_), .ZN(G1342gat));
  AOI21_X1  g688(.A(G134gat), .B1(new_n866_), .B2(new_n651_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n645_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(G134gat), .B2(new_n891_), .ZN(G1343gat));
  NAND3_X1  g691(.A1(new_n791_), .A2(new_n398_), .A3(new_n445_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT123), .Z(new_n894_));
  NOR2_X1   g693(.A1(new_n882_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n599_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n557_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT124), .B(G148gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1345gat));
  NAND2_X1  g699(.A1(new_n895_), .A2(new_n615_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  AOI21_X1  g702(.A(G162gat), .B1(new_n895_), .B2(new_n651_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n895_), .A2(G162gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n696_), .B2(new_n905_), .ZN(G1347gat));
  NOR3_X1   g705(.A1(new_n703_), .A2(new_n398_), .A3(new_n656_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n600_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n436_), .B(new_n909_), .C1(new_n841_), .C2(new_n854_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(G169gat), .A3(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n870_), .A2(new_n302_), .A3(new_n909_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n913_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n910_), .A2(G169gat), .A3(new_n916_), .A4(new_n911_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n915_), .A3(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n914_), .A2(new_n920_), .A3(new_n915_), .A4(new_n917_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1348gat));
  NAND2_X1  g721(.A1(new_n870_), .A2(new_n907_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n844_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n303_), .ZN(G1349gat));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n694_), .ZN(new_n926_));
  MUX2_X1   g725(.A(G183gat), .B(new_n276_), .S(new_n926_), .Z(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n923_), .B2(new_n645_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n651_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n923_), .B2(new_n929_), .ZN(G1351gat));
  NOR2_X1   g729(.A1(new_n882_), .A2(new_n455_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n656_), .A2(new_n397_), .A3(new_n436_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n600_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(new_n259_), .ZN(G1352gat));
  NOR2_X1   g734(.A1(new_n933_), .A2(new_n844_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(new_n257_), .ZN(G1353gat));
  INV_X1    g736(.A(new_n933_), .ZN(new_n938_));
  AOI211_X1 g737(.A(KEYINPUT63), .B(G211gat), .C1(new_n938_), .C2(new_n615_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT63), .B(G211gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n933_), .A2(new_n694_), .A3(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1354gat));
  XOR2_X1   g741(.A(KEYINPUT127), .B(G218gat), .Z(new_n943_));
  NOR3_X1   g742(.A1(new_n933_), .A2(new_n645_), .A3(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n938_), .A2(new_n651_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n943_), .ZN(G1355gat));
endmodule


