//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR3_X1   g004(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT66), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  OR3_X1    g006(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(new_n204_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n207_), .A2(new_n210_), .A3(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT8), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT10), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT10), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n220_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n229_));
  INV_X1    g028(.A(G85gat), .ZN(new_n230_));
  INV_X1    g029(.A(G92gat), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT9), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n215_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n208_), .A2(new_n204_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n218_), .B1(new_n235_), .B2(new_n215_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n219_), .A2(new_n234_), .A3(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(G57gat), .A2(G64gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G57gat), .A2(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G78gat), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n240_), .A2(new_n246_), .A3(new_n241_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n244_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n239_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n249_), .A2(new_n219_), .A3(new_n234_), .A4(new_n238_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(KEYINPUT12), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n239_), .A2(new_n250_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n203_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n202_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT5), .B(G176gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G204gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G120gat), .B(G148gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n253_), .A2(new_n255_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n202_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n257_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n263_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT67), .B1(new_n258_), .B2(new_n270_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n264_), .B(new_n266_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n272_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n258_), .A2(KEYINPUT67), .A3(new_n270_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n276_), .A2(new_n277_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(KEYINPUT13), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n275_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G15gat), .B(G22gat), .ZN(new_n282_));
  INV_X1    g081(.A(G1gat), .ZN(new_n283_));
  INV_X1    g082(.A(G8gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G1gat), .B(G8gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G29gat), .B(G36gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G43gat), .B(G50gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G43gat), .B(G50gat), .Z(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n289_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n288_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT15), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n295_), .B(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n296_), .B1(new_n298_), .B2(new_n288_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G229gat), .A2(G233gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n288_), .B(new_n295_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(G229gat), .A3(G233gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT75), .B(G169gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(G197gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G113gat), .B(G141gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n308_), .A2(KEYINPUT74), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n304_), .B(new_n309_), .Z(new_n310_));
  NAND2_X1  g109(.A1(new_n281_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT19), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT95), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT22), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(G169gat), .ZN(new_n319_));
  INV_X1    g118(.A(G169gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n320_), .A2(KEYINPUT22), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n317_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(KEYINPUT22), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(G169gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(KEYINPUT95), .ZN(new_n325_));
  AOI21_X1  g124(.A(G176gat), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G176gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n320_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT96), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT23), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G183gat), .A3(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n323_), .A2(new_n324_), .A3(KEYINPUT95), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT95), .B1(new_n323_), .B2(new_n324_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n327_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT96), .ZN(new_n341_));
  INV_X1    g140(.A(new_n328_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n329_), .A2(new_n337_), .A3(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT93), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT93), .ZN(new_n348_));
  AND2_X1   g147(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT26), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT94), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT24), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n328_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n357_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT94), .B1(new_n366_), .B2(new_n363_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n330_), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT79), .B1(new_n330_), .B2(KEYINPUT23), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n333_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(new_n361_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n365_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n344_), .A2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G197gat), .B(G204gat), .Z(new_n375_));
  INV_X1    g174(.A(KEYINPUT92), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G211gat), .A2(G218gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G211gat), .A2(G218gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n376_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(G211gat), .A2(G218gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(KEYINPUT92), .A3(new_n377_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n380_), .A2(new_n382_), .A3(KEYINPUT21), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT21), .B1(new_n380_), .B2(new_n382_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n375_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n382_), .A3(KEYINPUT21), .ZN(new_n386_));
  INV_X1    g185(.A(new_n375_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n316_), .B1(new_n374_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(new_n388_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n392_));
  INV_X1    g191(.A(new_n333_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n331_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n330_), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n393_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n392_), .B1(new_n397_), .B2(new_n335_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n399_));
  AOI21_X1  g198(.A(G176gat), .B1(new_n321_), .B2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n323_), .C1(new_n399_), .C2(new_n321_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n370_), .A2(KEYINPUT80), .A3(new_n336_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n398_), .A2(new_n401_), .A3(new_n342_), .A4(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n345_), .A2(new_n346_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n354_), .A2(KEYINPUT76), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n406_), .B(G190gat), .C1(new_n355_), .C2(KEYINPUT76), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT76), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n408_), .B(KEYINPUT26), .C1(new_n353_), .C2(KEYINPUT77), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n404_), .A2(new_n405_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n364_), .A2(new_n410_), .A3(new_n334_), .A4(new_n371_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n391_), .A2(new_n403_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n315_), .B1(new_n390_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n403_), .A2(new_n411_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n389_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n344_), .A2(new_n373_), .A3(new_n391_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n415_), .A2(KEYINPUT20), .A3(new_n315_), .A4(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT97), .B(KEYINPUT18), .Z(new_n419_));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n413_), .A2(new_n418_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n374_), .A2(new_n389_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(KEYINPUT20), .A3(new_n412_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n314_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n423_), .B1(new_n428_), .B2(new_n417_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n312_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT101), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT101), .B(new_n312_), .C1(new_n425_), .C2(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G127gat), .B(G134gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G113gat), .B(G120gat), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n439_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(KEYINPUT85), .A3(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n441_), .A2(KEYINPUT85), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G155gat), .ZN(new_n445_));
  INV_X1    g244(.A(G162gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(G141gat), .A2(G148gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(KEYINPUT3), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT3), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n453_), .B(KEYINPUT88), .C1(G141gat), .C2(G148gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT2), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n452_), .A2(new_n454_), .B1(KEYINPUT89), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G141gat), .A2(G148gat), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n457_), .A2(new_n455_), .A3(KEYINPUT89), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n459_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n449_), .B1(new_n456_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n450_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT1), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n447_), .A2(new_n465_), .A3(new_n448_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n448_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n467_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n464_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n444_), .B1(new_n462_), .B2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n462_), .A2(new_n469_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n440_), .A2(new_n441_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n437_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n462_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n464_), .A2(new_n468_), .A3(new_n466_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT4), .B1(new_n477_), .B2(new_n444_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n436_), .B1(new_n474_), .B2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n470_), .A2(new_n473_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n435_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G29gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G85gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT0), .B(G57gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n479_), .A2(new_n481_), .A3(new_n486_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT91), .B1(new_n493_), .B2(new_n391_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n389_), .B(new_n495_), .C1(new_n492_), .C2(new_n471_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G228gat), .A2(G233gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n497_), .B1(new_n471_), .B2(new_n492_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  NOR4_X1   g298(.A1(new_n462_), .A2(new_n469_), .A3(KEYINPUT29), .A4(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G78gat), .B(G106gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n498_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n475_), .A2(new_n492_), .A3(new_n476_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n499_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n471_), .A2(new_n492_), .A3(new_n497_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n501_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n494_), .B(new_n496_), .C1(new_n503_), .C2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n496_), .A2(new_n494_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n502_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G22gat), .B(G50gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  NAND3_X1  g314(.A1(new_n508_), .A2(new_n512_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n508_), .A2(new_n512_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n515_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT84), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n414_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n403_), .A2(new_n411_), .A3(new_n522_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n521_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G15gat), .B(G43gat), .ZN(new_n527_));
  AND2_X1   g326(.A1(G227gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G71gat), .B(G99gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n531_), .B(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n520_), .B1(new_n526_), .B2(new_n534_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n403_), .A2(new_n411_), .A3(new_n522_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n522_), .B1(new_n403_), .B2(new_n411_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT84), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n524_), .A2(new_n521_), .A3(new_n525_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n531_), .B(new_n532_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n444_), .B(KEYINPUT31), .Z(new_n542_));
  AND3_X1   g341(.A1(new_n535_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n535_), .B2(new_n541_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n516_), .B(new_n519_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n542_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT86), .B1(new_n538_), .B2(new_n540_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n535_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n508_), .A2(new_n515_), .A3(new_n512_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n515_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n549_), .B(new_n550_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n545_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT100), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n390_), .A2(new_n315_), .A3(new_n412_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n416_), .A2(KEYINPUT20), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT99), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT99), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n416_), .A2(new_n559_), .A3(KEYINPUT20), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n560_), .A3(new_n415_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n556_), .B1(new_n561_), .B2(new_n314_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n555_), .B1(new_n562_), .B2(new_n423_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n557_), .A2(KEYINPUT99), .B1(new_n414_), .B2(new_n389_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n315_), .B1(new_n564_), .B2(new_n560_), .ZN(new_n565_));
  OAI211_X1 g364(.A(KEYINPUT100), .B(new_n424_), .C1(new_n565_), .C2(new_n556_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n428_), .A2(new_n423_), .A3(new_n417_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n563_), .A2(KEYINPUT27), .A3(new_n566_), .A4(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n434_), .A2(new_n491_), .A3(new_n554_), .A4(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n489_), .A2(KEYINPUT33), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n479_), .A2(new_n481_), .A3(new_n571_), .A4(new_n486_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n424_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n435_), .B1(new_n474_), .B2(new_n478_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n486_), .B1(new_n480_), .B2(new_n436_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n573_), .A2(new_n567_), .A3(new_n574_), .A4(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n423_), .A2(KEYINPUT32), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n490_), .B1(new_n562_), .B2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n428_), .A2(new_n417_), .A3(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT98), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n428_), .A2(new_n583_), .A3(new_n417_), .A4(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n578_), .B1(new_n580_), .B2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n543_), .A2(new_n544_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n551_), .A2(new_n552_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n311_), .B1(new_n569_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n288_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(new_n250_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT72), .B(KEYINPUT16), .Z(new_n594_));
  XNOR2_X1  g393(.A(G127gat), .B(G155gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT17), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n593_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n593_), .B1(new_n601_), .B2(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT73), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606_));
  INV_X1    g405(.A(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT69), .B(G190gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT36), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT35), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n239_), .A2(new_n295_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT70), .B1(new_n298_), .B2(new_n239_), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n612_), .B(new_n615_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n615_), .A2(new_n612_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(new_n612_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n616_), .A2(new_n617_), .A3(new_n620_), .A4(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n611_), .B1(new_n618_), .B2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n616_), .A2(new_n617_), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n619_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n610_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n628_), .A3(new_n622_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(KEYINPUT71), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT37), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n624_), .A2(KEYINPUT71), .A3(KEYINPUT37), .A4(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n605_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n590_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n283_), .A3(new_n490_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT38), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n281_), .A2(new_n639_), .A3(new_n310_), .A4(new_n603_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n624_), .A2(new_n629_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n603_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT102), .B1(new_n311_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n569_), .A2(new_n589_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n491_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n638_), .A2(new_n648_), .ZN(G1324gat));
  XNOR2_X1  g448(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n434_), .A2(new_n568_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n643_), .A2(new_n645_), .A3(new_n652_), .A4(new_n646_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n654_), .A3(G8gat), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n653_), .A2(KEYINPUT104), .A3(new_n654_), .A4(G8gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n660_));
  AOI211_X1 g459(.A(new_n660_), .B(new_n654_), .C1(new_n653_), .C2(G8gat), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n653_), .A2(G8gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT103), .B1(new_n662_), .B2(KEYINPUT39), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n659_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n636_), .A2(new_n284_), .A3(new_n652_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n651_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n663_), .A2(new_n661_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n665_), .B(new_n650_), .C1(new_n668_), .C2(new_n659_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n647_), .B2(new_n587_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n587_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n636_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n676_), .ZN(G1326gat));
  INV_X1    g476(.A(G22gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n588_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n636_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n647_), .A2(new_n588_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(G22gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G22gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT107), .ZN(G1327gat));
  NOR2_X1   g485(.A1(new_n311_), .A2(new_n604_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n634_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n634_), .B2(new_n690_), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n688_), .B(new_n691_), .C1(new_n569_), .C2(new_n589_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n691_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n646_), .B2(new_n634_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n687_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(G29gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n491_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n687_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n646_), .A2(new_n634_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n691_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n646_), .A2(new_n634_), .A3(new_n693_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n698_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(KEYINPUT44), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n687_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT109), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n695_), .B(new_n697_), .C1(new_n704_), .C2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n604_), .A2(new_n642_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n590_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n696_), .B1(new_n711_), .B2(new_n491_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT110), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n708_), .A2(new_n715_), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1328gat));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n710_), .A2(new_n718_), .A3(new_n652_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT45), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n695_), .A2(new_n652_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n703_), .B1(new_n702_), .B2(KEYINPUT44), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n705_), .A2(KEYINPUT109), .A3(new_n706_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n724_), .B2(new_n718_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n720_), .B(KEYINPUT46), .C1(new_n724_), .C2(new_n718_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1329gat));
  INV_X1    g528(.A(G43gat), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n587_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n695_), .B(new_n731_), .C1(new_n704_), .C2(new_n707_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n711_), .B2(new_n587_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT47), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(new_n736_), .A3(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1330gat));
  AOI21_X1  g537(.A(G50gat), .B1(new_n710_), .B2(new_n679_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n695_), .ZN(new_n740_));
  AOI211_X1 g539(.A(new_n588_), .B(new_n740_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(G50gat), .ZN(G1331gat));
  INV_X1    g541(.A(new_n281_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n310_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n569_), .B2(new_n589_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n635_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n490_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(new_n642_), .A3(new_n604_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n751_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n490_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n749_), .B1(new_n754_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n748_), .A2(new_n756_), .A3(new_n652_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n752_), .A2(new_n652_), .A3(new_n753_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(G64gat), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G64gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1333gat));
  OR3_X1    g561(.A1(new_n747_), .A2(G71gat), .A3(new_n587_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n752_), .A2(new_n675_), .A3(new_n753_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G71gat), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(KEYINPUT49), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(KEYINPUT49), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1334gat));
  OR3_X1    g567(.A1(new_n747_), .A2(G78gat), .A3(new_n588_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n752_), .A2(new_n679_), .A3(new_n753_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(G78gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G78gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1335gat));
  INV_X1    g573(.A(new_n745_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n605_), .B(new_n775_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n491_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n746_), .A2(new_n709_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n230_), .A3(new_n490_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT113), .ZN(G1336gat));
  AOI21_X1  g580(.A(G92gat), .B1(new_n778_), .B2(new_n652_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n776_), .B1(new_n568_), .B2(new_n434_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(G92gat), .ZN(G1337gat));
  NAND2_X1  g583(.A1(new_n746_), .A2(new_n709_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n226_), .A2(new_n227_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(new_n587_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G99gat), .B1(new_n776_), .B2(new_n587_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT114), .B(G99gat), .C1(new_n776_), .C2(new_n587_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n793_), .B(new_n787_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1338gat));
  OAI21_X1  g596(.A(G106gat), .B1(new_n776_), .B2(new_n588_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n746_), .A2(new_n220_), .A3(new_n679_), .A4(new_n709_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT116), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT52), .B(G106gat), .C1(new_n776_), .C2(new_n588_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g604(.A1(new_n652_), .A2(new_n491_), .A3(new_n545_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n268_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT117), .B1(new_n256_), .B2(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n256_), .A2(KEYINPUT55), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n253_), .A2(new_n203_), .A3(new_n255_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .A4(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n263_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n276_), .A2(new_n277_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(new_n817_), .A3(new_n263_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n815_), .A2(new_n310_), .A3(new_n816_), .A4(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n278_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n299_), .A2(new_n300_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n302_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n300_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n308_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n304_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n308_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n819_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n642_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(KEYINPUT118), .A3(new_n642_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n818_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n817_), .B1(new_n813_), .B2(new_n263_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n837_), .A2(KEYINPUT58), .A3(new_n816_), .A4(new_n826_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n815_), .A2(new_n816_), .A3(new_n826_), .A4(new_n818_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n841_), .A3(new_n634_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n828_), .A2(KEYINPUT57), .A3(new_n642_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n603_), .B1(new_n834_), .B2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n635_), .A2(new_n744_), .A3(new_n281_), .ZN(new_n846_));
  XOR2_X1   g645(.A(new_n846_), .B(KEYINPUT54), .Z(new_n847_));
  OAI21_X1  g646(.A(new_n806_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT59), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT118), .B1(new_n828_), .B2(new_n642_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n830_), .B(new_n641_), .C1(new_n819_), .C2(new_n827_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n832_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n842_), .A2(new_n843_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n605_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n847_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n652_), .A2(KEYINPUT59), .A3(new_n491_), .A4(new_n545_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n849_), .A2(G113gat), .A3(new_n310_), .A4(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n310_), .B(new_n806_), .C1(new_n845_), .C2(new_n847_), .ZN(new_n861_));
  INV_X1    g660(.A(G113gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT120), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n861_), .A2(new_n865_), .A3(new_n862_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n860_), .A2(new_n864_), .A3(new_n866_), .ZN(G1340gat));
  NAND3_X1  g666(.A1(new_n849_), .A2(new_n743_), .A3(new_n859_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G120gat), .ZN(new_n869_));
  INV_X1    g668(.A(new_n848_), .ZN(new_n870_));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n281_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n870_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n871_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n869_), .A2(new_n873_), .ZN(G1341gat));
  NAND4_X1  g673(.A1(new_n849_), .A2(G127gat), .A3(new_n603_), .A4(new_n859_), .ZN(new_n875_));
  INV_X1    g674(.A(G127gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n848_), .B2(new_n605_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1342gat));
  INV_X1    g677(.A(G134gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n848_), .B2(new_n642_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT121), .B(new_n879_), .C1(new_n848_), .C2(new_n642_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n848_), .A2(KEYINPUT59), .B1(new_n857_), .B2(new_n858_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n634_), .A2(G134gat), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT122), .Z(new_n886_));
  AOI22_X1  g685(.A1(new_n882_), .A2(new_n883_), .B1(new_n884_), .B2(new_n886_), .ZN(G1343gat));
  NOR2_X1   g686(.A1(new_n652_), .A2(new_n491_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n553_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n644_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n856_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n310_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT123), .B(G141gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1344gat));
  NAND2_X1  g694(.A1(new_n892_), .A2(new_n743_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G148gat), .ZN(G1345gat));
  XOR2_X1   g696(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n445_), .B1(new_n892_), .B2(new_n604_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n890_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n604_), .B(new_n901_), .C1(new_n845_), .C2(new_n847_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(G155gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n899_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n892_), .A2(new_n445_), .A3(new_n604_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(G155gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(new_n906_), .A3(new_n898_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(G1346gat));
  AOI21_X1  g707(.A(G162gat), .B1(new_n892_), .B2(new_n641_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n845_), .A2(new_n847_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n910_), .A2(new_n688_), .A3(new_n890_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(G162gat), .B2(new_n911_), .ZN(G1347gat));
  AOI21_X1  g711(.A(new_n490_), .B1(new_n434_), .B2(new_n568_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n675_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n679_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n604_), .B1(new_n834_), .B2(new_n844_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n310_), .B(new_n915_), .C1(new_n916_), .C2(new_n847_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n338_), .A2(new_n339_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT62), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(G169gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n920_), .ZN(G1348gat));
  INV_X1    g722(.A(new_n915_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G176gat), .B1(new_n925_), .B2(new_n743_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n913_), .A2(new_n743_), .A3(new_n675_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n910_), .B2(new_n679_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n891_), .A2(new_n856_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n930_), .A2(KEYINPUT125), .A3(new_n588_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n927_), .B1(new_n929_), .B2(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n926_), .B1(new_n932_), .B2(G176gat), .ZN(G1349gat));
  AND4_X1   g732(.A1(new_n603_), .A2(new_n925_), .A3(new_n351_), .A4(new_n347_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n914_), .A2(new_n605_), .ZN(new_n935_));
  AOI21_X1  g734(.A(KEYINPUT125), .B1(new_n930_), .B2(new_n588_), .ZN(new_n936_));
  AOI211_X1 g735(.A(new_n928_), .B(new_n679_), .C1(new_n891_), .C2(new_n856_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(G183gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n934_), .B1(new_n938_), .B2(new_n939_), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n857_), .A2(new_n634_), .A3(new_n915_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(G190gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n641_), .A2(new_n358_), .ZN(new_n943_));
  AOI211_X1 g742(.A(new_n924_), .B(new_n943_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n945_), .A3(KEYINPUT126), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n353_), .B1(new_n925_), .B2(new_n634_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n944_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n946_), .A2(new_n949_), .ZN(G1351gat));
  AND2_X1   g749(.A1(new_n913_), .A2(new_n889_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n930_), .A2(new_n310_), .A3(new_n951_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g752(.A1(new_n930_), .A2(new_n743_), .A3(new_n951_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n930_), .A2(new_n603_), .A3(new_n951_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(KEYINPUT63), .B(G211gat), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n958_), .B1(new_n956_), .B2(new_n959_), .ZN(G1354gat));
  OAI211_X1 g759(.A(new_n641_), .B(new_n951_), .C1(new_n845_), .C2(new_n847_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(KEYINPUT127), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n930_), .A2(new_n963_), .A3(new_n641_), .A4(new_n951_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n962_), .A2(new_n964_), .A3(new_n607_), .ZN(new_n965_));
  NAND4_X1  g764(.A1(new_n930_), .A2(G218gat), .A3(new_n634_), .A4(new_n951_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1355gat));
endmodule


