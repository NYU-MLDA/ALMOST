//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT83), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT25), .B(G183gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT82), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT82), .B1(new_n219_), .B2(new_n220_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n210_), .B(new_n218_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(KEYINPUT84), .A2(G176gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT84), .A2(G176gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT22), .B(G169gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT85), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n228_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n204_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n215_), .A2(new_n232_), .A3(new_n216_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT86), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n223_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G99gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n235_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G113gat), .B(G120gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n238_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  INV_X1    g042(.A(G15gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT30), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT31), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n242_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT102), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n239_), .B(new_n240_), .Z(new_n253_));
  OR2_X1    g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT2), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT89), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n259_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265_));
  INV_X1    g064(.A(G141gat), .ZN(new_n266_));
  INV_X1    g065(.A(G148gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT88), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT88), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n265_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n256_), .B1(new_n264_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT87), .B1(new_n255_), .B2(KEYINPUT1), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT87), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(G155gat), .A4(G162gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n255_), .A2(KEYINPUT1), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n275_), .A2(new_n278_), .A3(new_n279_), .A4(new_n254_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n270_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n281_), .A2(new_n261_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n253_), .B1(new_n274_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n256_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n261_), .A2(new_n262_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT2), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n258_), .A2(new_n259_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n257_), .ZN(new_n289_));
  NOR4_X1   g088(.A1(KEYINPUT88), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n271_), .B1(new_n270_), .B2(new_n265_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n285_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n280_), .A2(new_n282_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(new_n241_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n284_), .A2(new_n295_), .A3(KEYINPUT101), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n274_), .A2(new_n283_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT101), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(new_n241_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(KEYINPUT4), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n284_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n252_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(new_n299_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT103), .B1(new_n304_), .B2(new_n252_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT103), .ZN(new_n306_));
  AOI211_X1 g105(.A(new_n306_), .B(new_n251_), .C1(new_n296_), .C2(new_n299_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n303_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G29gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(G85gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT0), .B(G57gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n300_), .A2(new_n302_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n251_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n304_), .A2(new_n252_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n306_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n304_), .A2(KEYINPUT103), .A3(new_n252_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n312_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n249_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G22gat), .B(G50gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327_));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G211gat), .B(G218gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT91), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G204gat), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n333_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n334_));
  INV_X1    g133(.A(G197gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(G204gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT21), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT90), .B1(new_n333_), .B2(G197gat), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n333_), .A2(G197gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT21), .B1(new_n341_), .B2(new_n336_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n332_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n334_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n329_), .A2(new_n344_), .A3(KEYINPUT21), .A4(new_n331_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n297_), .B2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(G228gat), .A2(G233gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n348_), .B1(KEYINPUT92), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G78gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G106gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n350_), .B(G78gat), .ZN(new_n354_));
  INV_X1    g153(.A(G106gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n326_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n297_), .A2(new_n347_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT28), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n349_), .A2(KEYINPUT92), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n353_), .A2(new_n356_), .A3(new_n326_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n362_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(new_n366_), .B2(new_n357_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n235_), .A2(new_n346_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT20), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n226_), .A2(new_n227_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n376_), .A2(KEYINPUT98), .A3(new_n204_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT98), .B1(new_n376_), .B2(new_n204_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n233_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n202_), .A2(KEYINPUT96), .A3(KEYINPUT24), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n380_), .A2(new_n207_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n202_), .A2(KEYINPUT24), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT96), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n217_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT95), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n220_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT26), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(G190gat), .ZN(new_n389_));
  INV_X1    g188(.A(G190gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(KEYINPUT26), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT95), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(new_n392_), .A3(new_n219_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n385_), .A2(KEYINPUT97), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT97), .B1(new_n385_), .B2(new_n393_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n379_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n375_), .B1(new_n346_), .B2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G8gat), .B(G36gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT99), .ZN(new_n404_));
  INV_X1    g203(.A(new_n374_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT20), .B1(new_n235_), .B2(new_n346_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT94), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n406_), .A2(new_n407_), .B1(new_n396_), .B2(new_n346_), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT94), .B(KEYINPUT20), .C1(new_n235_), .C2(new_n346_), .ZN(new_n409_));
  AOI211_X1 g208(.A(new_n404_), .B(new_n405_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n396_), .A2(new_n346_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT99), .B1(new_n413_), .B2(new_n374_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n397_), .B(new_n403_), .C1(new_n410_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT108), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n379_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n393_), .B2(new_n385_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n374_), .B1(new_n419_), .B2(new_n371_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(new_n413_), .B2(new_n374_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n415_), .A2(new_n416_), .B1(new_n402_), .B2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n369_), .B1(new_n417_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n397_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n402_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n369_), .A3(new_n415_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n368_), .B1(new_n423_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT109), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n368_), .B(KEYINPUT109), .C1(new_n423_), .C2(new_n427_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n324_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT33), .B1(new_n308_), .B2(new_n313_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n313_), .A2(KEYINPUT33), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n316_), .A2(new_n318_), .A3(new_n319_), .A4(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT104), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n296_), .A2(new_n436_), .A3(new_n299_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n251_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n315_), .A2(new_n252_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n312_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n433_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(new_n425_), .A3(new_n415_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT105), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n443_), .A2(new_n425_), .A3(KEYINPUT105), .A4(new_n415_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n403_), .A2(KEYINPUT32), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n397_), .B(new_n448_), .C1(new_n410_), .C2(new_n414_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n421_), .A2(KEYINPUT32), .A3(new_n403_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n322_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT106), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT106), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n322_), .A2(new_n453_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n446_), .A2(new_n447_), .A3(new_n452_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n368_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT107), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT107), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n458_), .A3(new_n368_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n423_), .A2(new_n427_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n322_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n364_), .A2(new_n367_), .A3(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n459_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n432_), .B1(new_n464_), .B2(new_n249_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G1gat), .A2(G8gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT14), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n468_), .B2(KEYINPUT75), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(KEYINPUT75), .B2(new_n468_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G1gat), .B(G8gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n470_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G29gat), .B(G36gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G43gat), .B(G50gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n473_), .B(new_n476_), .Z(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(G229gat), .A3(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT79), .ZN(new_n479_));
  INV_X1    g278(.A(new_n473_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n476_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n476_), .B(KEYINPUT15), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n473_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n484_), .B(KEYINPUT80), .Z(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G113gat), .B(G141gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT81), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G169gat), .B(G197gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  OR2_X1    g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n465_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n498_));
  XOR2_X1   g297(.A(G71gat), .B(G78gat), .Z(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n499_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(G231gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT76), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(new_n473_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G127gat), .B(G155gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G183gat), .B(G211gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT17), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(KEYINPUT78), .ZN(new_n515_));
  INV_X1    g314(.A(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(KEYINPUT17), .A3(new_n516_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT6), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n523_));
  OR3_X1    g322(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G85gat), .B(G92gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT64), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n526_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT64), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n525_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT8), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(KEYINPUT9), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT10), .B(G99gat), .Z(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n355_), .ZN(new_n535_));
  INV_X1    g334(.A(G85gat), .ZN(new_n536_));
  INV_X1    g335(.A(G92gat), .ZN(new_n537_));
  OR3_X1    g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT9), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n533_), .A2(new_n535_), .A3(new_n522_), .A4(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n532_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n503_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT12), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n540_), .A2(new_n503_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G230gat), .A2(G233gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n543_), .A2(KEYINPUT65), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n547_), .B2(new_n541_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n541_), .B2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G120gat), .B(G148gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G176gat), .B(G204gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT67), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n555_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n546_), .A2(new_n558_), .A3(new_n549_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n557_), .B(new_n559_), .C1(KEYINPUT68), .C2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n540_), .A2(new_n476_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT34), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n532_), .A2(new_n539_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n569_), .A2(KEYINPUT70), .A3(new_n482_), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT70), .B1(new_n569_), .B2(new_n482_), .ZN(new_n571_));
  OAI221_X1 g370(.A(new_n566_), .B1(KEYINPUT35), .B2(new_n568_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(KEYINPUT35), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT69), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n572_), .B(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G190gat), .B(G218gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT71), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT72), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n575_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n574_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n572_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n579_), .B(new_n580_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT73), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(new_n588_), .A3(KEYINPUT37), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT74), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n575_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(KEYINPUT74), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n593_), .A3(new_n587_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n583_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n590_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n496_), .A2(new_n520_), .A3(new_n565_), .A4(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n598_), .A2(G1gat), .A3(new_n461_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT38), .Z(new_n600_));
  INV_X1    g399(.A(new_n595_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n465_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n565_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n520_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n495_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT110), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(KEYINPUT110), .A3(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G1gat), .B1(new_n611_), .B2(new_n461_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n600_), .A2(new_n612_), .ZN(G1324gat));
  INV_X1    g412(.A(new_n460_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G8gat), .B1(new_n606_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT39), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n598_), .A2(G8gat), .A3(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(KEYINPUT40), .A3(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1325gat));
  INV_X1    g421(.A(KEYINPUT111), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT41), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n610_), .A2(new_n248_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(G15gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n249_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n627_), .A2(KEYINPUT41), .A3(new_n244_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n623_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n624_), .A3(G15gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT41), .B1(new_n627_), .B2(new_n244_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(KEYINPUT111), .A3(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n598_), .A2(G15gat), .A3(new_n249_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT112), .Z(new_n634_));
  NAND3_X1  g433(.A1(new_n629_), .A2(new_n632_), .A3(new_n634_), .ZN(G1326gat));
  OR3_X1    g434(.A1(new_n598_), .A2(G22gat), .A3(new_n368_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G22gat), .B1(new_n611_), .B2(new_n368_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT42), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT42), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n636_), .B1(new_n638_), .B2(new_n639_), .ZN(G1327gat));
  NAND2_X1  g439(.A1(new_n601_), .A2(new_n604_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n603_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n496_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n322_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT43), .B1(new_n465_), .B2(new_n597_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  INV_X1    g445(.A(new_n597_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n458_), .B1(new_n455_), .B2(new_n368_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n460_), .A2(new_n462_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n248_), .B1(new_n650_), .B2(new_n459_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n646_), .B(new_n647_), .C1(new_n651_), .C2(new_n432_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n645_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n565_), .A2(new_n604_), .A3(new_n494_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT44), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n657_), .B(new_n654_), .C1(new_n645_), .C2(new_n652_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n322_), .A2(G29gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n644_), .B1(new_n659_), .B2(new_n660_), .ZN(G1328gat));
  XNOR2_X1  g460(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n656_), .A2(new_n658_), .A3(new_n614_), .ZN(new_n664_));
  INV_X1    g463(.A(G36gat), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND4_X1   g465(.A1(new_n665_), .A2(new_n496_), .A3(new_n460_), .A4(new_n642_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT45), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n663_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n668_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n670_), .B(new_n662_), .C1(new_n665_), .C2(new_n664_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1329gat));
  AOI21_X1  g471(.A(G43gat), .B1(new_n643_), .B2(new_n248_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n248_), .A2(G43gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n659_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT47), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(G1330gat));
  INV_X1    g476(.A(G50gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n368_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n643_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT114), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n659_), .A2(new_n681_), .A3(new_n679_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G50gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n659_), .B2(new_n679_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1331gat));
  NOR2_X1   g484(.A1(new_n465_), .A2(new_n494_), .ZN(new_n686_));
  AND4_X1   g485(.A1(new_n520_), .A2(new_n686_), .A3(new_n603_), .A4(new_n597_), .ZN(new_n687_));
  INV_X1    g486(.A(G57gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n322_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n602_), .A2(new_n520_), .A3(new_n495_), .A4(new_n603_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n461_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1332gat));
  OAI21_X1  g491(.A(G64gat), .B1(new_n690_), .B2(new_n614_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT48), .ZN(new_n694_));
  INV_X1    g493(.A(G64gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n695_), .A3(new_n460_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1333gat));
  OAI21_X1  g496(.A(G71gat), .B1(new_n690_), .B2(new_n249_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT49), .ZN(new_n699_));
  INV_X1    g498(.A(G71gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n687_), .A2(new_n700_), .A3(new_n248_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1334gat));
  OAI21_X1  g501(.A(G78gat), .B1(new_n690_), .B2(new_n368_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT50), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n687_), .A2(new_n351_), .A3(new_n679_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1335gat));
  NAND3_X1  g505(.A1(new_n603_), .A2(new_n604_), .A3(new_n495_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n653_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n461_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n641_), .A2(new_n565_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n686_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n322_), .A2(new_n536_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(G1336gat));
  OAI21_X1  g513(.A(G92gat), .B1(new_n709_), .B2(new_n614_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n460_), .A2(new_n537_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n712_), .B2(new_n716_), .ZN(G1337gat));
  OAI21_X1  g516(.A(G99gat), .B1(new_n709_), .B2(new_n249_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n248_), .A2(new_n534_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g520(.A(new_n432_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n455_), .A2(new_n458_), .A3(new_n368_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n723_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(new_n248_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n646_), .B1(new_n725_), .B2(new_n647_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n465_), .A2(KEYINPUT43), .A3(new_n597_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n679_), .B(new_n708_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT116), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n653_), .A2(KEYINPUT116), .A3(new_n679_), .A4(new_n708_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n730_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n731_), .ZN(new_n732_));
  AND4_X1   g531(.A1(new_n355_), .A2(new_n686_), .A3(new_n679_), .A4(new_n711_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT115), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n368_), .B(new_n707_), .C1(new_n645_), .C2(new_n652_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n355_), .B1(new_n736_), .B2(KEYINPUT116), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT52), .B1(new_n737_), .B2(new_n730_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT53), .B1(new_n735_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  INV_X1    g539(.A(new_n730_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n731_), .A2(G106gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n732_), .A4(new_n734_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n739_), .A2(new_n745_), .ZN(G1339gat));
  NAND2_X1  g545(.A1(new_n494_), .A2(new_n559_), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n544_), .A2(KEYINPUT118), .A3(new_n545_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n546_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n544_), .A2(KEYINPUT55), .A3(new_n545_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT118), .B1(new_n544_), .B2(new_n545_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n748_), .A2(new_n750_), .A3(new_n751_), .A4(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n556_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(KEYINPUT119), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(KEYINPUT119), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n753_), .A2(new_n556_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n747_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n477_), .A2(new_n485_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n485_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n481_), .A2(new_n483_), .A3(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n491_), .A3(new_n762_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n560_), .A2(new_n492_), .A3(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n595_), .B1(new_n759_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT120), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n754_), .A2(new_n768_), .A3(KEYINPUT56), .ZN(new_n769_));
  XNOR2_X1  g568(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n753_), .A2(new_n556_), .A3(new_n770_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n492_), .A2(new_n559_), .A3(new_n763_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n769_), .A2(KEYINPUT58), .A3(new_n771_), .A4(new_n772_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n647_), .A3(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT57), .B(new_n595_), .C1(new_n759_), .C2(new_n764_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n767_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n604_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n495_), .A2(new_n781_), .A3(new_n520_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT117), .B1(new_n604_), .B2(new_n494_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n597_), .A2(new_n782_), .A3(new_n565_), .A4(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n780_), .A2(new_n787_), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n461_), .B(new_n249_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT59), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n495_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(G113gat), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(KEYINPUT121), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n790_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n494_), .A2(new_n796_), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n795_), .A2(new_n796_), .B1(new_n800_), .B2(new_n801_), .ZN(G1340gat));
  AOI21_X1  g601(.A(new_n565_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n803_));
  INV_X1    g602(.A(G120gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n565_), .B2(KEYINPUT60), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(KEYINPUT60), .B2(new_n804_), .ZN(new_n806_));
  OAI22_X1  g605(.A1(new_n803_), .A2(new_n804_), .B1(new_n800_), .B2(new_n806_), .ZN(G1341gat));
  AOI21_X1  g606(.A(new_n604_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n808_));
  INV_X1    g607(.A(G127gat), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n520_), .A2(new_n809_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n808_), .A2(new_n809_), .B1(new_n800_), .B2(new_n810_), .ZN(G1342gat));
  NAND3_X1  g610(.A1(new_n797_), .A2(new_n601_), .A3(new_n799_), .ZN(new_n812_));
  INV_X1    g611(.A(G134gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n792_), .A2(new_n794_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n647_), .A2(G134gat), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT122), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n812_), .A2(new_n813_), .B1(new_n814_), .B2(new_n816_), .ZN(G1343gat));
  NAND4_X1  g616(.A1(new_n614_), .A2(new_n322_), .A3(new_n249_), .A4(new_n679_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT123), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n788_), .A2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(new_n495_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(new_n266_), .ZN(G1344gat));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n565_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(new_n267_), .ZN(G1345gat));
  AND2_X1   g623(.A1(new_n788_), .A2(new_n819_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT124), .A3(new_n520_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n820_), .B2(new_n604_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT61), .B(G155gat), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n826_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1346gat));
  OR3_X1    g631(.A1(new_n820_), .A2(G162gat), .A3(new_n595_), .ZN(new_n833_));
  OAI21_X1  g632(.A(G162gat), .B1(new_n820_), .B2(new_n597_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(G1347gat));
  NOR3_X1   g634(.A1(new_n614_), .A2(new_n679_), .A3(new_n324_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n788_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT126), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n786_), .B1(new_n779_), .B2(new_n604_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n836_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT126), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n838_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n227_), .A3(new_n494_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n839_), .A2(new_n495_), .A3(new_n840_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n205_), .B1(new_n846_), .B2(KEYINPUT125), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT125), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n837_), .B2(new_n495_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n847_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n845_), .B1(new_n851_), .B2(new_n852_), .ZN(G1348gat));
  NOR3_X1   g652(.A1(new_n837_), .A2(new_n206_), .A3(new_n565_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n844_), .A2(new_n603_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n226_), .ZN(G1349gat));
  AOI21_X1  g655(.A(G183gat), .B1(new_n841_), .B2(new_n520_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n604_), .A2(new_n219_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n844_), .B2(new_n858_), .ZN(G1350gat));
  INV_X1    g658(.A(new_n844_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n601_), .A2(new_n392_), .A3(new_n387_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n597_), .B1(new_n838_), .B2(new_n843_), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n860_), .A2(new_n861_), .B1(new_n862_), .B2(new_n390_), .ZN(G1351gat));
  NOR3_X1   g662(.A1(new_n614_), .A2(new_n248_), .A3(new_n462_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n788_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n495_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(new_n335_), .ZN(G1352gat));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n565_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n333_), .ZN(G1353gat));
  AND2_X1   g668(.A1(new_n788_), .A2(new_n864_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n520_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n872_));
  AND2_X1   g671(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n871_), .B2(new_n872_), .ZN(G1354gat));
  OR3_X1    g674(.A1(new_n865_), .A2(G218gat), .A3(new_n595_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G218gat), .B1(new_n865_), .B2(new_n597_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1355gat));
endmodule


