//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n204_));
  OR2_X1    g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT84), .ZN(new_n209_));
  OR2_X1    g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(KEYINPUT1), .B2(new_n207_), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n205_), .B(new_n206_), .C1(new_n209_), .C2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT85), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT85), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n205_), .A2(KEYINPUT86), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT3), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n206_), .A2(KEYINPUT87), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n218_), .B(KEYINPUT2), .Z(new_n219_));
  AOI22_X1  g018(.A1(new_n217_), .A2(new_n219_), .B1(G155gat), .B2(G162gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n210_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G127gat), .B(G134gat), .Z(new_n223_));
  XOR2_X1   g022(.A(G113gat), .B(G120gat), .Z(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT83), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n224_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n223_), .A2(new_n224_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n215_), .A2(new_n226_), .A3(new_n229_), .A4(new_n221_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n204_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n215_), .A2(new_n221_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT93), .B(KEYINPUT4), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n232_), .A2(new_n227_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n203_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n228_), .A2(new_n230_), .A3(new_n202_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT0), .B(G57gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G85gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(G1gat), .B(G29gat), .Z(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT33), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G226gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT19), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT20), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT26), .B(G190gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT79), .ZN(new_n250_));
  INV_X1    g049(.A(G183gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(KEYINPUT25), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT25), .B(G183gat), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n249_), .B(new_n252_), .C1(new_n253_), .C2(new_n250_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT80), .ZN(new_n255_));
  INV_X1    g054(.A(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT24), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT81), .Z(new_n262_));
  MUX2_X1   g061(.A(new_n262_), .B(new_n261_), .S(KEYINPUT23), .Z(new_n263_));
  OR2_X1    g062(.A1(new_n258_), .A2(KEYINPUT24), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n255_), .A2(new_n260_), .A3(new_n263_), .A4(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n262_), .B2(KEYINPUT23), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n267_), .B1(G183gat), .B2(G190gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n259_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT22), .B(G169gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(new_n257_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n265_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(G197gat), .B(G204gat), .Z(new_n275_));
  OAI21_X1  g074(.A(new_n274_), .B1(new_n275_), .B2(KEYINPUT21), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT21), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n248_), .B1(new_n273_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n263_), .B1(G183gat), .B2(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT92), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n271_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n249_), .A2(new_n253_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n260_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n286_), .A2(KEYINPUT90), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(KEYINPUT90), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n287_), .A2(new_n267_), .A3(new_n264_), .A4(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT91), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n247_), .B(new_n280_), .C1(new_n291_), .C2(new_n279_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT18), .B(G64gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(G92gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n279_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT20), .B1(new_n273_), .B2(new_n279_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT89), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n299_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n297_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n292_), .B(new_n296_), .C1(new_n303_), .C2(new_n247_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n292_), .B1(new_n303_), .B2(new_n247_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n296_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n228_), .A2(new_n230_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n242_), .B1(new_n308_), .B2(new_n203_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n231_), .A2(new_n234_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n310_), .B2(new_n203_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n244_), .A2(new_n304_), .A3(new_n307_), .A4(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n296_), .A2(KEYINPUT32), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT94), .Z(new_n314_));
  OAI211_X1 g113(.A(new_n292_), .B(new_n314_), .C1(new_n303_), .C2(new_n247_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n284_), .A2(new_n278_), .A3(new_n289_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n280_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n246_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(new_n302_), .B2(new_n246_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n313_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n235_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n243_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n315_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT95), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT95), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n315_), .A2(new_n320_), .A3(new_n325_), .A4(new_n322_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n312_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G78gat), .B(G106gat), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n278_), .B1(new_n222_), .B2(KEYINPUT29), .ZN(new_n330_));
  INV_X1    g129(.A(G228gat), .ZN(new_n331_));
  INV_X1    g130(.A(G233gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n330_), .A2(new_n334_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n329_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT88), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT28), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n341_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n337_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n335_), .A3(new_n328_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n338_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n227_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n273_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G71gat), .B(G99gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT31), .ZN(new_n355_));
  XOR2_X1   g154(.A(G15gat), .B(G43gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G227gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n353_), .B(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n338_), .A2(new_n347_), .A3(KEYINPUT88), .A4(new_n344_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n349_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n353_), .B(new_n359_), .Z(new_n364_));
  AOI22_X1  g163(.A1(new_n340_), .A2(new_n344_), .B1(new_n347_), .B2(new_n338_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n361_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n322_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n367_), .A2(new_n362_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT27), .B1(new_n307_), .B2(new_n304_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n319_), .A2(new_n306_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n304_), .A2(new_n371_), .A3(KEYINPUT27), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n327_), .A2(new_n363_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G15gat), .B(G22gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT75), .B(G8gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT14), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G1gat), .ZN(new_n379_));
  INV_X1    g178(.A(G1gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(new_n377_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G8gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G29gat), .ZN(new_n385_));
  INV_X1    g184(.A(G36gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G43gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G29gat), .A2(G36gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G50gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n388_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G29gat), .B(G36gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G43gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(G50gat), .B1(new_n396_), .B2(new_n390_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n384_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n382_), .B(G8gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n398_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G229gat), .A3(G233gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n392_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n396_), .A2(G50gat), .A3(new_n390_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n405_), .A2(KEYINPUT15), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT15), .B1(new_n405_), .B2(new_n406_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n400_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G229gat), .A2(G233gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n399_), .A3(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G113gat), .B(G141gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(new_n256_), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(G197gat), .Z(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n404_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n404_), .B2(new_n412_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT13), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G85gat), .A2(G92gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT65), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT9), .ZN(new_n424_));
  INV_X1    g223(.A(G85gat), .ZN(new_n425_));
  INV_X1    g224(.A(G92gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT9), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n421_), .A2(new_n422_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431_));
  INV_X1    g230(.A(G99gat), .ZN(new_n432_));
  INV_X1    g231(.A(G106gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(KEYINPUT10), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT10), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G99gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n433_), .A2(KEYINPUT64), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT64), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n430_), .A2(new_n436_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT66), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT67), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n434_), .A2(new_n453_), .A3(new_n435_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n448_), .A2(new_n455_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n427_), .A2(new_n421_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n446_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G64gat), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n465_));
  XOR2_X1   g264(.A(G71gat), .B(G78gat), .Z(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n465_), .A2(new_n466_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n462_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n446_), .B(new_n469_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT68), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G230gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n457_), .A2(new_n459_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT8), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT68), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n446_), .A4(new_n469_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n475_), .A3(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n483_));
  NAND2_X1  g282(.A1(new_n471_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT69), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n446_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n430_), .A2(KEYINPUT69), .A3(new_n436_), .A4(new_n445_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(KEYINPUT12), .A3(new_n470_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n484_), .A2(new_n474_), .A3(new_n472_), .A4(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G120gat), .B(G148gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(G176gat), .B(G204gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  AND3_X1   g295(.A1(new_n482_), .A2(new_n491_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n482_), .B2(new_n491_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n420_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n482_), .A2(new_n491_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n482_), .A2(new_n491_), .A3(new_n496_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(KEYINPUT13), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT74), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n506_), .A2(KEYINPUT37), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(KEYINPUT37), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G232gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT34), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n407_), .A2(new_n408_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n479_), .B2(new_n488_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n398_), .B(new_n446_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OAI211_X1 g313(.A(KEYINPUT35), .B(new_n510_), .C1(new_n512_), .C2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n489_), .A2(new_n409_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(KEYINPUT35), .ZN(new_n517_));
  INV_X1    g316(.A(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n516_), .A2(new_n517_), .A3(new_n520_), .A4(new_n513_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT72), .B(G134gat), .ZN(new_n522_));
  INV_X1    g321(.A(G162gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G190gat), .B(G218gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n527_));
  AND4_X1   g326(.A1(new_n515_), .A2(new_n521_), .A3(new_n526_), .A4(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n526_), .B(KEYINPUT36), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n515_), .B2(new_n521_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n507_), .B(new_n508_), .C1(new_n528_), .C2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n400_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n400_), .A2(new_n533_), .ZN(new_n535_));
  OR3_X1    g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n470_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n470_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G127gat), .B(G155gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n540_), .B(new_n541_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n544_), .A2(KEYINPUT17), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n536_), .A2(new_n537_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551_));
  INV_X1    g350(.A(new_n547_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n545_), .A2(new_n546_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n548_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  AOI211_X1 g356(.A(new_n519_), .B(new_n518_), .C1(new_n516_), .C2(new_n513_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n521_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n529_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n515_), .A2(new_n521_), .A3(new_n526_), .A4(new_n527_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n560_), .A2(new_n506_), .A3(KEYINPUT37), .A4(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n532_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  NOR4_X1   g362(.A1(new_n374_), .A2(new_n419_), .A3(new_n505_), .A4(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n322_), .B(KEYINPUT96), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n380_), .A3(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT38), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n528_), .A2(new_n531_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT98), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n374_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n557_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n505_), .A2(new_n419_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT97), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n573_), .A2(new_n368_), .A3(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n568_), .B1(new_n380_), .B2(new_n576_), .ZN(G1324gat));
  INV_X1    g376(.A(new_n557_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n374_), .A2(new_n578_), .A3(new_n571_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n575_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n373_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n579_), .A2(KEYINPUT99), .A3(new_n580_), .A4(new_n581_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(G8gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT39), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n584_), .A2(new_n585_), .A3(new_n588_), .A4(G8gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n376_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n564_), .A2(new_n591_), .A3(new_n581_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT40), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(KEYINPUT40), .A3(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(G1325gat));
  INV_X1    g396(.A(G15gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n564_), .A2(new_n598_), .A3(new_n364_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n573_), .A2(new_n575_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n364_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n601_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT41), .B1(new_n601_), .B2(G15gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT100), .B(new_n599_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1326gat));
  INV_X1    g407(.A(G22gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n349_), .A2(new_n361_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n600_), .B2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT42), .Z(new_n612_));
  NAND3_X1  g411(.A1(new_n564_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(G1327gat));
  NAND2_X1  g413(.A1(new_n327_), .A2(new_n363_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n369_), .A2(new_n373_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT43), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n532_), .A2(new_n562_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT43), .B1(new_n374_), .B2(new_n619_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n580_), .A3(new_n578_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT44), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n623_), .A2(KEYINPUT44), .A3(new_n580_), .A4(new_n578_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n566_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT101), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n626_), .A2(new_n630_), .A3(new_n566_), .A4(new_n627_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(G29gat), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n569_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n557_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n617_), .A2(new_n574_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT102), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n617_), .A2(new_n637_), .A3(new_n574_), .A4(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n385_), .A3(new_n322_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n632_), .A2(new_n641_), .ZN(G1328gat));
  NAND3_X1  g441(.A1(new_n626_), .A2(new_n581_), .A3(new_n627_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G36gat), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n636_), .A2(new_n386_), .A3(new_n581_), .A4(new_n638_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT45), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n644_), .A2(KEYINPUT46), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1329gat));
  NAND3_X1  g450(.A1(new_n626_), .A2(new_n364_), .A3(new_n627_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G43gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n640_), .A2(new_n388_), .A3(new_n364_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT47), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(KEYINPUT47), .A3(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1330gat));
  NAND3_X1  g458(.A1(new_n640_), .A2(new_n392_), .A3(new_n610_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n626_), .A2(new_n610_), .A3(new_n627_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(new_n392_), .ZN(G1331gat));
  INV_X1    g461(.A(new_n505_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n617_), .A2(new_n664_), .A3(new_n419_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n419_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT103), .B1(new_n374_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n663_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n532_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G57gat), .B1(new_n670_), .B2(new_n566_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n663_), .A2(new_n666_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n573_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n368_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n671_), .B1(G57gat), .B2(new_n676_), .ZN(G1332gat));
  INV_X1    g476(.A(G64gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n670_), .A2(new_n678_), .A3(new_n581_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n581_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G64gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT104), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n683_), .A3(G64gat), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n682_), .A2(KEYINPUT48), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT48), .B1(new_n682_), .B2(new_n684_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n679_), .B1(new_n685_), .B2(new_n686_), .ZN(G1333gat));
  INV_X1    g486(.A(G71gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n670_), .A2(new_n688_), .A3(new_n364_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT49), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n674_), .A2(new_n364_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(G71gat), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT49), .B(new_n688_), .C1(new_n674_), .C2(new_n364_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(G1334gat));
  INV_X1    g495(.A(G78gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n670_), .A2(new_n697_), .A3(new_n610_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n610_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G78gat), .B1(new_n675_), .B2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(KEYINPUT50), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(KEYINPUT50), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(G1335gat));
  NAND2_X1  g502(.A1(new_n668_), .A2(new_n634_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT106), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n668_), .A2(new_n706_), .A3(new_n634_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G85gat), .B1(new_n708_), .B2(new_n566_), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n557_), .B(new_n673_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(new_n322_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(G85gat), .B2(new_n711_), .ZN(G1336gat));
  NAND3_X1  g511(.A1(new_n708_), .A2(new_n426_), .A3(new_n581_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n710_), .A2(new_n581_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n713_), .B(new_n714_), .C1(new_n426_), .C2(new_n715_), .ZN(new_n716_));
  AOI211_X1 g515(.A(G92gat), .B(new_n373_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(new_n426_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT107), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1337gat));
  NAND3_X1  g519(.A1(new_n708_), .A2(new_n440_), .A3(new_n364_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n710_), .A2(new_n364_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n721_), .B(new_n722_), .C1(new_n432_), .C2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n440_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n725_), .B(new_n360_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n723_), .A2(new_n432_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT51), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n724_), .A2(new_n728_), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n708_), .A2(new_n444_), .A3(new_n610_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT53), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n623_), .A2(new_n578_), .A3(new_n610_), .A4(new_n672_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G106gat), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n733_), .A2(new_n732_), .A3(G106gat), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n730_), .B(new_n731_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n444_), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n737_), .B(new_n699_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n735_), .A2(new_n734_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT53), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(new_n740_), .ZN(G1339gat));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n610_), .A2(new_n360_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AND4_X1   g543(.A1(G229gat), .A2(new_n410_), .A3(new_n399_), .A4(G233gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n411_), .B2(new_n403_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n417_), .B1(new_n415_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n490_), .A2(new_n472_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n483_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n462_), .B2(new_n470_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n475_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n491_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n491_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT55), .A3(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT56), .B1(new_n756_), .B2(new_n501_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n758_), .B(new_n496_), .C1(new_n753_), .C2(new_n755_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n503_), .B(new_n747_), .C1(new_n757_), .C2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT113), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n619_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n484_), .A2(new_n472_), .A3(new_n490_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n475_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n754_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n765_), .A2(new_n764_), .A3(new_n475_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n501_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n758_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n496_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT56), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n497_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(KEYINPUT58), .A4(new_n747_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n762_), .A2(new_n763_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n747_), .B1(new_n498_), .B2(new_n497_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT112), .B1(new_n778_), .B2(KEYINPUT56), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n501_), .B(new_n779_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(KEYINPUT112), .A2(KEYINPUT56), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n666_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n503_), .B1(new_n771_), .B2(new_n779_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n777_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n633_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n784_), .A2(KEYINPUT57), .A3(new_n633_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n776_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n578_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n499_), .A2(new_n504_), .A3(new_n419_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n669_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT109), .B1(new_n792_), .B2(KEYINPUT54), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n499_), .A2(new_n504_), .A3(new_n419_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT109), .B(KEYINPUT54), .C1(new_n794_), .C2(new_n563_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n563_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT108), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n794_), .A2(new_n563_), .A3(new_n800_), .A4(KEYINPUT54), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n793_), .A2(new_n796_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n795_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(KEYINPUT110), .C1(new_n799_), .C2(new_n801_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n744_), .B1(new_n790_), .B2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n581_), .A2(new_n565_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT59), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n789_), .A2(new_n578_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  INV_X1    g613(.A(new_n811_), .ZN(new_n815_));
  NOR4_X1   g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .A4(new_n744_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n742_), .B1(new_n812_), .B2(new_n816_), .ZN(new_n817_));
  OR2_X1    g616(.A1(KEYINPUT115), .A2(G113gat), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n804_), .A2(new_n808_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n784_), .A2(KEYINPUT57), .A3(new_n633_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT57), .B1(new_n784_), .B2(new_n633_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n557_), .B1(new_n822_), .B2(new_n776_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n811_), .B(new_n743_), .C1(new_n819_), .C2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n814_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n810_), .A2(KEYINPUT59), .A3(new_n811_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(KEYINPUT114), .ZN(new_n827_));
  OAI21_X1  g626(.A(G113gat), .B1(new_n419_), .B2(KEYINPUT115), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n817_), .A2(new_n818_), .A3(new_n827_), .A4(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(G113gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n824_), .B2(new_n419_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT116), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n834_), .A3(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1340gat));
  INV_X1    g635(.A(new_n824_), .ZN(new_n837_));
  INV_X1    g636(.A(G120gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n663_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n837_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n838_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n663_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n838_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n837_), .B2(new_n557_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n817_), .A2(new_n827_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n557_), .A2(G127gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g647(.A(G134gat), .B1(new_n837_), .B2(new_n571_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT118), .B(G134gat), .Z(new_n850_));
  NOR2_X1   g649(.A1(new_n619_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n846_), .B2(new_n851_), .ZN(G1343gat));
  NOR3_X1   g651(.A1(new_n813_), .A2(new_n699_), .A3(new_n364_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n811_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n666_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g656(.A1(new_n854_), .A2(new_n663_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT119), .B(G148gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1345gat));
  NOR2_X1   g659(.A1(new_n854_), .A2(new_n578_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT61), .B(G155gat), .Z(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT120), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n861_), .B(new_n863_), .ZN(G1346gat));
  NOR3_X1   g663(.A1(new_n854_), .A2(new_n523_), .A3(new_n619_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n855_), .A2(new_n571_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n523_), .B2(new_n866_), .ZN(G1347gat));
  NOR3_X1   g666(.A1(new_n813_), .A2(new_n566_), .A3(new_n744_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n581_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT121), .A3(new_n666_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n869_), .B2(new_n419_), .ZN(new_n873_));
  AND2_X1   g672(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n871_), .A2(G169gat), .A3(new_n873_), .A4(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n666_), .A2(new_n270_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT123), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n870_), .A2(new_n877_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n871_), .A2(G169gat), .A3(new_n873_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n875_), .B(new_n878_), .C1(new_n879_), .C2(new_n880_), .ZN(G1348gat));
  AND2_X1   g680(.A1(KEYINPUT124), .A2(G176gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(KEYINPUT124), .A2(G176gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n869_), .A2(new_n663_), .ZN(new_n885_));
  MUX2_X1   g684(.A(new_n882_), .B(new_n884_), .S(new_n885_), .Z(G1349gat));
  NOR2_X1   g685(.A1(new_n869_), .A2(new_n578_), .ZN(new_n887_));
  MUX2_X1   g686(.A(G183gat), .B(new_n253_), .S(new_n887_), .Z(G1350gat));
  NAND3_X1  g687(.A1(new_n870_), .A2(new_n571_), .A3(new_n249_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n870_), .A2(new_n620_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n890_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT125), .B1(new_n890_), .B2(G190gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n889_), .B1(new_n891_), .B2(new_n892_), .ZN(G1351gat));
  NOR2_X1   g692(.A1(new_n373_), .A2(new_n322_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n853_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n666_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n505_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n896_), .B(new_n557_), .C1(new_n901_), .C2(new_n902_), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n895_), .A2(new_n578_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT126), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n903_), .A2(new_n907_), .A3(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1354gat));
  AOI21_X1  g708(.A(G218gat), .B1(new_n896_), .B2(new_n571_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n620_), .A2(G218gat), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT127), .Z(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n896_), .B2(new_n912_), .ZN(G1355gat));
endmodule


