//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G71gat), .ZN(new_n205_));
  INV_X1    g004(.A(G78gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT69), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n202_), .A2(new_n203_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n209_), .A2(KEYINPUT69), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(KEYINPUT69), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(new_n211_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT68), .ZN(new_n218_));
  XOR2_X1   g017(.A(G85gat), .B(G92gat), .Z(new_n219_));
  AND2_X1   g018(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n221_));
  OAI22_X1  g020(.A1(new_n220_), .A2(new_n221_), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(KEYINPUT67), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT6), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT67), .B1(new_n222_), .B2(new_n226_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n219_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n222_), .A2(new_n232_), .A3(new_n226_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n219_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT66), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n236_), .A2(new_n240_), .A3(new_n237_), .A4(new_n219_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(KEYINPUT8), .A2(new_n235_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n243_));
  XOR2_X1   g042(.A(KEYINPUT10), .B(G99gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n225_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT64), .B(G92gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT9), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(G85gat), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n243_), .A2(new_n245_), .A3(new_n232_), .A4(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n218_), .B1(new_n242_), .B2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n239_), .A2(new_n241_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n222_), .A2(new_n226_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(new_n232_), .A3(new_n227_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n237_), .B1(new_n256_), .B2(new_n219_), .ZN(new_n257_));
  OAI211_X1 g056(.A(KEYINPUT68), .B(new_n249_), .C1(new_n252_), .C2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n217_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n213_), .A2(new_n216_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT70), .B1(new_n252_), .B2(new_n257_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n242_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n260_), .B1(new_n264_), .B2(new_n249_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n259_), .B1(new_n265_), .B2(KEYINPUT12), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G230gat), .A2(G233gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n251_), .A2(new_n217_), .A3(new_n258_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT71), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n268_), .A2(KEYINPUT71), .A3(new_n269_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n266_), .B(new_n267_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n259_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n268_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n267_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G120gat), .B(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT5), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G176gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G204gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n281_), .B(KEYINPUT72), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n277_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT13), .ZN(new_n287_));
  INV_X1    g086(.A(G228gat), .ZN(new_n288_));
  INV_X1    g087(.A(G233gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n293_), .B(new_n294_), .C1(new_n297_), .C2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n295_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n294_), .B(KEYINPUT1), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n303_), .B(new_n298_), .C1(new_n304_), .C2(new_n292_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT29), .ZN(new_n307_));
  INV_X1    g106(.A(G204gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT91), .ZN(new_n310_));
  INV_X1    g109(.A(G197gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(G204gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(G204gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n309_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G211gat), .B(G218gat), .Z(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT21), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT92), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(KEYINPUT90), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n308_), .A2(G197gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(new_n311_), .B2(G204gat), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n318_), .B(KEYINPUT21), .C1(new_n319_), .C2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT21), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n323_), .B(new_n309_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n315_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n314_), .A2(new_n327_), .A3(KEYINPUT21), .A4(new_n315_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n317_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n291_), .B1(new_n307_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT94), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT93), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n317_), .A2(KEYINPUT93), .A3(new_n326_), .A4(new_n328_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AND4_X1   g135(.A1(new_n332_), .A2(new_n336_), .A3(new_n291_), .A4(new_n307_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n290_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(new_n338_), .B2(new_n307_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n331_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G78gat), .B(G106gat), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G22gat), .B(G50gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  OR3_X1    g144(.A1(new_n306_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT89), .B1(new_n306_), .B2(KEYINPUT29), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n349_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n345_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n346_), .A2(new_n347_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n348_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(new_n344_), .A3(new_n350_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n341_), .B(new_n331_), .C1(new_n337_), .C2(new_n339_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n343_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT97), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n343_), .A2(new_n357_), .A3(KEYINPUT97), .A4(new_n358_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT86), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n365_), .A2(KEYINPUT23), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(KEYINPUT23), .ZN(new_n367_));
  OAI22_X1  g166(.A1(new_n366_), .A2(new_n367_), .B1(G183gat), .B2(G190gat), .ZN(new_n368_));
  INV_X1    g167(.A(G176gat), .ZN(new_n369_));
  AND2_X1   g168(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT82), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT22), .B(G169gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n369_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n368_), .A2(new_n373_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n381_));
  OAI211_X1 g180(.A(KEYINPUT24), .B(new_n377_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT25), .B(G183gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT26), .B(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT24), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(new_n379_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n365_), .B(KEYINPUT23), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n382_), .A2(new_n385_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n378_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n378_), .B2(new_n392_), .ZN(new_n395_));
  INV_X1    g194(.A(G227gat), .ZN(new_n396_));
  OAI22_X1  g195(.A1(new_n394_), .A2(new_n395_), .B1(new_n396_), .B2(new_n289_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n378_), .A2(new_n392_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT85), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n396_), .A2(new_n289_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n378_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G15gat), .B(G43gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT84), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G71gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n397_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G99gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n407_), .A2(new_n408_), .A3(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n400_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n405_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n397_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n410_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n364_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G120gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G127gat), .B(G134gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G113gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n420_), .A2(G113gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(G120gat), .A3(new_n421_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(KEYINPUT31), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n411_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n415_), .A2(new_n410_), .A3(new_n416_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(KEYINPUT86), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n418_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n427_), .A2(new_n306_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n424_), .A2(new_n426_), .A3(new_n305_), .A4(new_n301_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(KEYINPUT102), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT102), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n427_), .A2(new_n440_), .A3(new_n306_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n436_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n437_), .A2(KEYINPUT4), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n435_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n439_), .A2(new_n441_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n434_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(G85gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT0), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G57gat), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n444_), .A2(new_n446_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n364_), .B(new_n428_), .C1(new_n412_), .C2(new_n417_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n433_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n336_), .A2(new_n291_), .A3(new_n307_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT94), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n338_), .A2(new_n332_), .A3(new_n307_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n330_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT96), .B1(new_n459_), .B2(new_n341_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT95), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n358_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT96), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n340_), .A2(new_n463_), .A3(new_n342_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n457_), .A2(new_n458_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n465_), .A2(KEYINPUT95), .A3(new_n341_), .A4(new_n331_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n460_), .A2(new_n462_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n357_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT18), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(G64gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n472_), .B(G92gat), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT19), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n372_), .A2(new_n377_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT100), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT100), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n372_), .A2(new_n481_), .A3(new_n377_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n368_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT101), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n480_), .A2(KEYINPUT101), .A3(new_n368_), .A4(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n377_), .A2(KEYINPUT24), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n488_), .A2(KEYINPUT98), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(KEYINPUT98), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n489_), .B(new_n490_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n386_), .A2(new_n389_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n391_), .A2(KEYINPUT99), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT99), .B1(new_n391_), .B2(new_n492_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n385_), .B(new_n491_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n487_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n478_), .B1(new_n496_), .B2(new_n329_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n398_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n334_), .A2(new_n498_), .A3(new_n335_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n477_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n329_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n487_), .A2(new_n501_), .A3(new_n495_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(KEYINPUT20), .A3(new_n477_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n498_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n474_), .B1(new_n500_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n494_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n391_), .A2(KEYINPUT99), .A3(new_n492_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n507_), .A2(new_n508_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n491_), .A2(new_n509_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT20), .B1(new_n510_), .B2(new_n501_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n499_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n476_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n336_), .A2(new_n398_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n514_), .A2(KEYINPUT20), .A3(new_n477_), .A4(new_n502_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n473_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT27), .B1(new_n506_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n495_), .A2(new_n483_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT20), .B1(new_n518_), .B2(new_n329_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT104), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT104), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n521_), .B(KEYINPUT20), .C1(new_n518_), .C2(new_n329_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n514_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n476_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n497_), .A2(new_n477_), .A3(new_n499_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n473_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n500_), .A2(new_n505_), .A3(new_n474_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n517_), .B1(new_n528_), .B2(KEYINPUT27), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n363_), .A2(new_n455_), .A3(new_n469_), .A4(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT106), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n363_), .A2(new_n469_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n453_), .A3(new_n529_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT105), .ZN(new_n535_));
  INV_X1    g334(.A(new_n453_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n473_), .A2(KEYINPUT32), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n513_), .A2(new_n537_), .A3(new_n515_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT103), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n538_), .A2(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n524_), .A2(new_n525_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(new_n537_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n452_), .B(KEYINPUT33), .ZN(new_n545_));
  OR3_X1    g344(.A1(new_n442_), .A2(new_n435_), .A3(new_n443_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n546_), .B(new_n450_), .C1(new_n434_), .C2(new_n445_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(new_n516_), .A3(new_n506_), .ZN(new_n548_));
  OAI22_X1  g347(.A1(new_n542_), .A2(new_n544_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n361_), .A2(new_n362_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(KEYINPUT27), .B(new_n516_), .C1(new_n543_), .C2(new_n473_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n517_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n363_), .B2(new_n469_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT105), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n453_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n535_), .A2(new_n551_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n433_), .A2(new_n454_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n532_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G29gat), .B(G36gat), .ZN(new_n561_));
  INV_X1    g360(.A(G43gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(G50gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n561_), .B(G43gat), .ZN(new_n565_));
  INV_X1    g364(.A(G50gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G1gat), .B(G8gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT76), .ZN(new_n572_));
  INV_X1    g371(.A(G15gat), .ZN(new_n573_));
  INV_X1    g372(.A(G22gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G15gat), .A2(G22gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G1gat), .A2(G8gat), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n575_), .A2(new_n576_), .B1(KEYINPUT14), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n572_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n570_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT79), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n568_), .B(KEYINPUT15), .Z(new_n583_));
  INV_X1    g382(.A(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n570_), .A2(new_n579_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n581_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n586_), .B1(new_n588_), .B2(new_n582_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G113gat), .B(G141gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(G169gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n311_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n586_), .B(new_n594_), .C1(new_n588_), .C2(new_n582_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(KEYINPUT80), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n595_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT80), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AOI211_X1 g398(.A(new_n287_), .B(new_n560_), .C1(new_n596_), .C2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n264_), .A2(new_n249_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n583_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n251_), .A2(new_n258_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT73), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT34), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(KEYINPUT35), .A3(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT74), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(G134gat), .ZN(new_n612_));
  INV_X1    g411(.A(G162gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT36), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n608_), .A2(KEYINPUT35), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n608_), .A2(KEYINPUT35), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n602_), .A2(new_n617_), .A3(new_n618_), .A4(new_n604_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n609_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT75), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n609_), .A2(KEYINPUT75), .A3(new_n616_), .A4(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n609_), .A2(new_n619_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n614_), .B(KEYINPUT36), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(KEYINPUT37), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n624_), .B2(new_n627_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n579_), .B(new_n633_), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(new_n260_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT16), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(G183gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(G211gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT17), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n635_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT77), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n639_), .A2(KEYINPUT17), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n635_), .A2(new_n640_), .A3(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n632_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n600_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT107), .ZN(new_n649_));
  INV_X1    g448(.A(G1gat), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n536_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT38), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n628_), .B(KEYINPUT108), .Z(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n560_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n287_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n597_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n645_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n453_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n651_), .A2(KEYINPUT38), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n652_), .A2(new_n660_), .A3(new_n661_), .ZN(G1324gat));
  OAI21_X1  g461(.A(KEYINPUT109), .B1(new_n659_), .B2(new_n529_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n657_), .A2(new_n654_), .A3(new_n560_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT109), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n664_), .A2(new_n665_), .A3(new_n645_), .A4(new_n554_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(G8gat), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT39), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n663_), .A2(new_n669_), .A3(G8gat), .A4(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G8gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n649_), .A2(new_n672_), .A3(new_n554_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n671_), .A2(new_n673_), .A3(KEYINPUT40), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1325gat));
  INV_X1    g477(.A(new_n559_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n649_), .A2(new_n573_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G15gat), .B1(new_n659_), .B2(new_n559_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT110), .Z(new_n682_));
  AND2_X1   g481(.A1(new_n682_), .A2(KEYINPUT41), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(KEYINPUT41), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1326gat));
  NAND3_X1  g484(.A1(new_n649_), .A2(new_n574_), .A3(new_n533_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G22gat), .B1(new_n659_), .B2(new_n550_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT42), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n556_), .B1(new_n555_), .B2(new_n453_), .ZN(new_n691_));
  NOR4_X1   g490(.A1(new_n550_), .A2(KEYINPUT105), .A3(new_n554_), .A4(new_n536_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n679_), .B1(new_n693_), .B2(new_n551_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n690_), .B(new_n632_), .C1(new_n694_), .C2(new_n532_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n632_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n560_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n646_), .A3(new_n658_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n698_), .A2(KEYINPUT44), .A3(new_n646_), .A4(new_n658_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n536_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n704_), .A2(KEYINPUT111), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(KEYINPUT111), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(G29gat), .A3(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n645_), .A2(new_n628_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n600_), .A2(new_n708_), .ZN(new_n709_));
  OR3_X1    g508(.A1(new_n709_), .A2(G29gat), .A3(new_n453_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  AND4_X1   g511(.A1(new_n712_), .A2(new_n600_), .A3(new_n554_), .A4(new_n708_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n701_), .A2(new_n554_), .A3(new_n702_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(G36gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G36gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n715_), .B(KEYINPUT46), .C1(new_n718_), .C2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1329gat));
  NAND3_X1  g523(.A1(new_n703_), .A2(G43gat), .A3(new_n679_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n562_), .B1(new_n709_), .B2(new_n559_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g527(.A(new_n566_), .B1(new_n703_), .B2(new_n533_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n709_), .A2(G50gat), .A3(new_n550_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1331gat));
  INV_X1    g530(.A(new_n597_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n287_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n560_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(new_n647_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n453_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n737_), .B(new_n738_), .C1(new_n736_), .C2(new_n735_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n599_), .A2(new_n645_), .A3(new_n596_), .ZN(new_n740_));
  NOR4_X1   g539(.A1(new_n560_), .A2(new_n656_), .A3(new_n654_), .A4(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n453_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n739_), .A2(new_n743_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT114), .Z(G1332gat));
  INV_X1    g544(.A(G64gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n741_), .B2(new_n554_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT48), .Z(new_n748_));
  NAND3_X1  g547(.A1(new_n735_), .A2(new_n746_), .A3(new_n554_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1333gat));
  AOI21_X1  g549(.A(new_n205_), .B1(new_n741_), .B2(new_n679_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT49), .Z(new_n752_));
  NAND3_X1  g551(.A1(new_n735_), .A2(new_n205_), .A3(new_n679_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1334gat));
  AOI21_X1  g553(.A(new_n206_), .B1(new_n741_), .B2(new_n533_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n735_), .A2(new_n206_), .A3(new_n533_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1335gat));
  AND2_X1   g558(.A1(new_n734_), .A2(new_n708_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n536_), .ZN(new_n761_));
  AOI211_X1 g560(.A(new_n645_), .B(new_n733_), .C1(new_n695_), .C2(new_n697_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n536_), .A2(G85gat), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT116), .Z(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n762_), .B2(new_n764_), .ZN(G1336gat));
  AOI21_X1  g564(.A(G92gat), .B1(new_n760_), .B2(new_n554_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n554_), .A2(new_n246_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n762_), .B2(new_n767_), .ZN(G1337gat));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(KEYINPUT51), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(KEYINPUT51), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n760_), .A2(new_n244_), .A3(new_n679_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT117), .Z(new_n773_));
  NAND2_X1  g572(.A1(new_n762_), .A2(new_n679_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G99gat), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n770_), .B(new_n771_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n776_));
  AND4_X1   g575(.A1(new_n769_), .A2(new_n773_), .A3(KEYINPUT51), .A4(new_n775_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1338gat));
  NAND3_X1  g577(.A1(new_n760_), .A2(new_n225_), .A3(new_n533_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n733_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n698_), .A2(new_n646_), .A3(new_n533_), .A4(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G106gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n779_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT119), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(new_n779_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n786_), .A2(KEYINPUT53), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT53), .B1(new_n786_), .B2(new_n788_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1339gat));
  NAND2_X1  g590(.A1(new_n597_), .A2(new_n282_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n284_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n265_), .A2(KEYINPUT12), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n273_), .B(new_n795_), .C1(new_n271_), .C2(new_n270_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n796_), .B2(new_n275_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n272_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n268_), .A2(new_n269_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT71), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n268_), .A2(KEYINPUT71), .A3(new_n269_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n804_), .A2(KEYINPUT55), .A3(new_n267_), .A4(new_n266_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n793_), .B1(new_n799_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n267_), .B1(new_n804_), .B2(new_n266_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n272_), .B1(new_n811_), .B2(new_n794_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n284_), .B1(new_n812_), .B2(new_n805_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT121), .B1(new_n813_), .B2(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(KEYINPUT56), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n792_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n582_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n581_), .A2(new_n818_), .A3(new_n585_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n592_), .B(new_n819_), .C1(new_n588_), .C2(new_n818_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n595_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n286_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT57), .B(new_n628_), .C1(new_n817_), .C2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT123), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n815_), .A2(new_n816_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n792_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n822_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n628_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n282_), .A2(new_n595_), .A3(new_n820_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n807_), .A2(new_n809_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n816_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n632_), .B1(new_n833_), .B2(KEYINPUT58), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(KEYINPUT58), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n632_), .B(KEYINPUT122), .C1(new_n833_), .C2(KEYINPUT58), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n810_), .A2(new_n814_), .B1(KEYINPUT56), .B2(new_n813_), .ZN(new_n840_));
  OAI22_X1  g639(.A1(new_n840_), .A2(new_n792_), .B1(new_n286_), .B2(new_n821_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(KEYINPUT57), .A4(new_n628_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n824_), .A2(new_n830_), .A3(new_n839_), .A4(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n740_), .B(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n656_), .A3(new_n696_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT54), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n847_), .A2(KEYINPUT54), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n844_), .A2(new_n646_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n533_), .A2(new_n554_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n536_), .A3(new_n679_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853_), .B2(new_n597_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n844_), .A2(new_n646_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n849_), .A2(new_n848_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n852_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n856_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n850_), .A2(KEYINPUT59), .A3(new_n852_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n855_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n859_), .A2(new_n856_), .A3(new_n860_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT59), .B1(new_n850_), .B2(new_n852_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(KEYINPUT124), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n863_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(G113gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n599_), .B2(new_n596_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n854_), .B1(new_n867_), .B2(new_n869_), .ZN(G1340gat));
  OAI21_X1  g669(.A(new_n419_), .B1(new_n656_), .B2(KEYINPUT60), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n419_), .A2(KEYINPUT60), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(KEYINPUT125), .B2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n853_), .B(new_n873_), .C1(KEYINPUT125), .C2(new_n871_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n861_), .A2(new_n862_), .A3(new_n656_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n419_), .ZN(G1341gat));
  AOI21_X1  g675(.A(G127gat), .B1(new_n853_), .B2(new_n645_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n645_), .A2(G127gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n867_), .B2(new_n878_), .ZN(G1342gat));
  AOI21_X1  g678(.A(G134gat), .B1(new_n853_), .B2(new_n654_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n632_), .A2(G134gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n867_), .B2(new_n881_), .ZN(G1343gat));
  NOR2_X1   g681(.A1(new_n850_), .A2(new_n679_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n883_), .A2(new_n536_), .A3(new_n555_), .A4(new_n597_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g684(.A1(new_n883_), .A2(new_n536_), .A3(new_n555_), .A4(new_n287_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g686(.A1(new_n883_), .A2(new_n536_), .A3(new_n645_), .A4(new_n555_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1346gat));
  AND3_X1   g689(.A1(new_n883_), .A2(new_n536_), .A3(new_n555_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n654_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n696_), .A2(new_n613_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n892_), .A2(new_n613_), .B1(new_n891_), .B2(new_n893_), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n850_), .A2(new_n533_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n529_), .A2(new_n536_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n559_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n895_), .A2(new_n374_), .A3(new_n597_), .A4(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n597_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT126), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n895_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n902_), .A2(new_n903_), .A3(G169gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n902_), .B2(G169gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n899_), .B1(new_n904_), .B2(new_n905_), .ZN(G1348gat));
  NAND3_X1  g705(.A1(new_n895_), .A2(new_n287_), .A3(new_n898_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g707(.A1(new_n895_), .A2(new_n645_), .A3(new_n898_), .ZN(new_n909_));
  MUX2_X1   g708(.A(new_n383_), .B(G183gat), .S(new_n909_), .Z(G1350gat));
  NAND2_X1  g709(.A1(new_n895_), .A2(new_n898_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G190gat), .B1(new_n911_), .B2(new_n696_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n654_), .A2(new_n384_), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT127), .Z(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n911_), .B2(new_n914_), .ZN(G1351gat));
  NOR3_X1   g714(.A1(new_n850_), .A2(new_n679_), .A3(new_n897_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n916_), .A2(new_n533_), .A3(new_n597_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n533_), .A3(new_n287_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n916_), .A2(new_n533_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n646_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT63), .B(G211gat), .Z(new_n924_));
  NAND4_X1  g723(.A1(new_n916_), .A2(new_n645_), .A3(new_n533_), .A4(new_n924_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1354gat));
  AND2_X1   g725(.A1(new_n916_), .A2(new_n533_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n654_), .ZN(new_n928_));
  INV_X1    g727(.A(G218gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n696_), .A2(new_n929_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n928_), .A2(new_n929_), .B1(new_n927_), .B2(new_n930_), .ZN(G1355gat));
endmodule


