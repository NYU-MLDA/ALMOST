//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  XOR2_X1   g007(.A(G29gat), .B(G36gat), .Z(new_n209_));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n211_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n206_), .B(new_n207_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT76), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n211_), .B(KEYINPUT15), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n214_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n212_), .A3(new_n219_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G113gat), .B(G141gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(G169gat), .B(G197gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n221_), .B(new_n224_), .C1(new_n229_), .C2(new_n228_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n236_));
  NOR2_X1   g035(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n238_), .A2(KEYINPUT80), .A3(new_n241_), .A4(new_n243_), .ZN(new_n248_));
  INV_X1    g047(.A(G176gat), .ZN(new_n249_));
  INV_X1    g048(.A(G169gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT79), .B1(new_n250_), .B2(KEYINPUT22), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT22), .B(G169gat), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n249_), .B(new_n251_), .C1(new_n252_), .C2(KEYINPUT79), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .A4(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G183gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT25), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G183gat), .ZN(new_n258_));
  INV_X1    g057(.A(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT26), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT26), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(G190gat), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n256_), .A2(new_n258_), .A3(new_n260_), .A4(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT24), .A3(new_n247_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT24), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n239_), .A2(KEYINPUT23), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(new_n239_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n254_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G15gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n274_), .B(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G127gat), .B(G134gat), .Z(new_n278_));
  XOR2_X1   g077(.A(G113gat), .B(G120gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n277_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G71gat), .B(G99gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT82), .B(G43gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n282_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT85), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT84), .B(KEYINPUT3), .ZN(new_n293_));
  INV_X1    g092(.A(G141gat), .ZN(new_n294_));
  INV_X1    g093(.A(G148gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n292_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT3), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n299_), .A2(KEYINPUT84), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(KEYINPUT84), .ZN(new_n301_));
  OAI211_X1 g100(.A(KEYINPUT85), .B(new_n298_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT2), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(G141gat), .A3(G148gat), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n304_), .A2(new_n306_), .B1(new_n296_), .B2(KEYINPUT3), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n297_), .A2(new_n302_), .A3(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n310_), .A2(KEYINPUT86), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT86), .B1(new_n310_), .B2(new_n311_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n296_), .A2(new_n303_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n309_), .B1(KEYINPUT1), .B2(new_n311_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n311_), .A2(KEYINPUT1), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT87), .B1(new_n315_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322_));
  AOI211_X1 g121(.A(new_n322_), .B(new_n319_), .C1(new_n308_), .C2(new_n314_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT28), .B1(new_n324_), .B2(KEYINPUT29), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n326_), .B(new_n327_), .C1(new_n321_), .C2(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT91), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n325_), .A2(new_n333_), .A3(new_n328_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G22gat), .B(G50gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT88), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n315_), .A2(new_n320_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n322_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n319_), .B1(new_n308_), .B2(new_n314_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT87), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(KEYINPUT29), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT21), .ZN(new_n345_));
  AND2_X1   g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT89), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(KEYINPUT89), .B(new_n345_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n346_), .A2(new_n347_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT21), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G211gat), .B(G218gat), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .A4(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n353_), .A2(new_n354_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT90), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT90), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n356_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n339_), .B1(new_n344_), .B2(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n355_), .A2(new_n356_), .ZN(new_n364_));
  AOI211_X1 g163(.A(new_n338_), .B(new_n364_), .C1(KEYINPUT29), .C2(new_n340_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n336_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n321_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n338_), .B1(new_n367_), .B2(new_n361_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n365_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n336_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n335_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n332_), .A2(new_n366_), .A3(new_n371_), .A4(new_n334_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G8gat), .B(G36gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT99), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n274_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n247_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n252_), .B2(new_n249_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(new_n272_), .B2(new_n242_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n238_), .A2(new_n241_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n364_), .B(new_n387_), .C1(new_n269_), .C2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n384_), .A2(KEYINPUT20), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n388_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT25), .B(G183gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT26), .B(G190gat), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n395_), .A2(new_n396_), .B1(new_n267_), .B2(new_n264_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT92), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n394_), .A2(new_n397_), .A3(new_n398_), .A4(new_n266_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT92), .B1(new_n269_), .B2(new_n388_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT93), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n387_), .A2(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(KEYINPUT93), .B(new_n386_), .C1(new_n272_), .C2(new_n242_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n357_), .B1(new_n401_), .B2(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n355_), .A2(new_n356_), .A3(new_n359_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n359_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n273_), .B(new_n254_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n392_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n406_), .A2(new_n409_), .A3(KEYINPUT20), .A4(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n383_), .B1(new_n393_), .B2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n411_), .A2(new_n383_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n382_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n254_), .A2(new_n273_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n361_), .B2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n410_), .B1(new_n417_), .B2(new_n406_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n399_), .A2(new_n400_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n419_), .A2(new_n364_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n384_), .A2(new_n420_), .A3(KEYINPUT20), .A4(new_n410_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n381_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n414_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n341_), .A2(new_n343_), .A3(new_n281_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(KEYINPUT4), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n315_), .A2(new_n320_), .A3(new_n280_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT95), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT95), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n342_), .A2(new_n433_), .A3(new_n280_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n324_), .A2(new_n281_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT96), .B1(new_n435_), .B2(KEYINPUT4), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n434_), .ZN(new_n437_));
  AND4_X1   g236(.A1(KEYINPUT96), .A2(new_n428_), .A3(new_n437_), .A4(KEYINPUT4), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n430_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n426_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G1gat), .B(G29gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G57gat), .B(G85gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  NAND3_X1  g244(.A1(new_n439_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n428_), .A2(new_n437_), .A3(KEYINPUT4), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT96), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n428_), .A2(new_n437_), .A3(KEYINPUT96), .A4(KEYINPUT4), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n429_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n440_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n447_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n425_), .B1(new_n446_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n446_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n447_), .A2(new_n456_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n439_), .A2(new_n440_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n380_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n406_), .A2(KEYINPUT20), .A3(new_n409_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n392_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n380_), .A3(new_n421_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n428_), .A2(KEYINPUT4), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(new_n427_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n445_), .B1(new_n435_), .B2(new_n427_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n465_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n457_), .A2(new_n459_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT98), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n455_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n457_), .A2(new_n470_), .A3(KEYINPUT98), .A4(new_n459_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n375_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n446_), .A2(new_n454_), .A3(new_n374_), .A4(new_n373_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT27), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n423_), .B2(new_n380_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n460_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n465_), .A2(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT100), .B1(new_n476_), .B2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n446_), .A2(new_n454_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT100), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n479_), .A2(new_n478_), .B1(new_n465_), .B2(new_n477_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n375_), .A4(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n291_), .B1(new_n475_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n375_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n486_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n290_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n234_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G57gat), .B(G64gat), .Z(new_n496_));
  INV_X1    g295(.A(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(KEYINPUT69), .B(G71gat), .Z(new_n499_));
  INV_X1    g298(.A(G78gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT69), .B(G71gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G78gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n498_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n504_), .A2(KEYINPUT70), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n496_), .A2(new_n497_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(KEYINPUT70), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT10), .B(G99gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(G106gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(G85gat), .B(G92gat), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT9), .ZN(new_n516_));
  INV_X1    g315(.A(G99gat), .ZN(new_n517_));
  INV_X1    g316(.A(G106gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT6), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT6), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(G99gat), .A3(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT9), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(G85gat), .A3(G92gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n516_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT72), .B1(new_n514_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT72), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n527_), .B(new_n528_), .C1(G106gat), .C2(new_n513_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT66), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n531_), .B(new_n532_), .C1(G99gat), .C2(G106gat), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n517_), .B(new_n518_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n522_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT8), .B1(new_n536_), .B2(new_n515_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n535_), .B(KEYINPUT68), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n522_), .B(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n515_), .A2(KEYINPUT8), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n537_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n530_), .B1(KEYINPUT71), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(KEYINPUT71), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT12), .B(new_n510_), .C1(new_n544_), .C2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT12), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n505_), .A2(new_n507_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n506_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n527_), .B1(G106gat), .B2(new_n513_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n543_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n548_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT64), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n555_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n547_), .A2(new_n556_), .A3(new_n558_), .A4(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n543_), .A2(new_n554_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n510_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n559_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n558_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT5), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G176gat), .B(G204gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n560_), .A2(new_n565_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT13), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n571_), .A2(KEYINPUT13), .A3(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n510_), .A2(new_n214_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n553_), .A2(new_n208_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n580_), .A2(new_n581_), .A3(G231gat), .A4(G233gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G127gat), .B(G155gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT16), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n586_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n590_), .A2(new_n591_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n585_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n580_), .A2(new_n581_), .B1(G231gat), .B2(G233gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT75), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n586_), .A2(new_n599_), .A3(new_n594_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n593_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT73), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT36), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT34), .ZN(new_n608_));
  OAI22_X1  g407(.A1(new_n561_), .A2(new_n213_), .B1(KEYINPUT35), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n541_), .A2(new_n542_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n537_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT71), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n545_), .A3(new_n530_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n609_), .B1(new_n615_), .B2(new_n222_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n608_), .A2(KEYINPUT35), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n616_), .A2(new_n618_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n606_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n621_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n605_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT36), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n619_), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n622_), .A2(new_n626_), .A3(KEYINPUT74), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT37), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n622_), .A2(new_n626_), .A3(KEYINPUT74), .A4(KEYINPUT37), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n495_), .A2(new_n579_), .A3(new_n601_), .A4(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n484_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n203_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n633_), .A2(KEYINPUT101), .A3(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT101), .B1(new_n633_), .B2(new_n635_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(KEYINPUT38), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n622_), .A2(new_n626_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n601_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n578_), .A2(new_n640_), .A3(new_n234_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n465_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n468_), .A2(new_n469_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n459_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n450_), .A2(new_n451_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n453_), .B1(new_n645_), .B2(new_n430_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT33), .B1(new_n646_), .B2(new_n445_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n472_), .B1(new_n644_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n454_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n452_), .A2(new_n453_), .A3(new_n447_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n414_), .B(new_n424_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n474_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n490_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n483_), .A2(new_n487_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n290_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n639_), .B(new_n641_), .C1(new_n655_), .C2(new_n493_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n488_), .B1(new_n490_), .B2(new_n652_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n494_), .B1(new_n659_), .B2(new_n290_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n660_), .A2(KEYINPUT102), .A3(new_n639_), .A4(new_n641_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n484_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n638_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT38), .B1(new_n636_), .B2(new_n637_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1324gat));
  OAI21_X1  g466(.A(G8gat), .B1(new_n656_), .B2(new_n486_), .ZN(new_n668_));
  XOR2_X1   g467(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n633_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n204_), .A3(new_n482_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n673_), .B(new_n675_), .ZN(G1325gat));
  INV_X1    g475(.A(G15gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n662_), .B2(new_n290_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT41), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n290_), .A2(new_n677_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n633_), .B2(new_n680_), .ZN(G1326gat));
  INV_X1    g480(.A(G22gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n375_), .A2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT106), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n671_), .A2(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n686_));
  INV_X1    g485(.A(new_n639_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT102), .B1(new_n688_), .B2(new_n641_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n656_), .A2(new_n657_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n375_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n686_), .B1(new_n691_), .B2(G22gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n490_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n686_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n693_), .A2(new_n682_), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n685_), .B1(new_n692_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT107), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n698_), .B(new_n685_), .C1(new_n692_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1327gat));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n629_), .A2(new_n702_), .A3(new_n630_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n655_), .B2(new_n493_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n631_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n706_), .A2(KEYINPUT43), .B1(new_n660_), .B2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n578_), .A2(new_n234_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n640_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n701_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n712_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n707_), .B1(new_n660_), .B2(new_n705_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n708_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT44), .B(new_n714_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n713_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G29gat), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n484_), .A2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n601_), .A2(new_n639_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(new_n578_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n495_), .A2(new_n634_), .A3(new_n723_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n718_), .A2(new_n720_), .B1(new_n719_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(KEYINPUT109), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n713_), .A2(new_n482_), .A3(new_n717_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G36gat), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n233_), .B(new_n723_), .C1(new_n655_), .C2(new_n493_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n486_), .A2(G36gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT45), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n495_), .A2(new_n735_), .A3(new_n723_), .A4(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n726_), .A2(KEYINPUT109), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n728_), .B1(new_n730_), .B2(new_n740_), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n727_), .B(new_n739_), .C1(new_n729_), .C2(G36gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1329gat));
  NAND4_X1  g542(.A1(new_n713_), .A2(G43gat), .A3(new_n717_), .A4(new_n290_), .ZN(new_n744_));
  INV_X1    g543(.A(G43gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n745_), .B1(new_n731_), .B2(new_n291_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n744_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g549(.A(G50gat), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n490_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n495_), .A2(new_n375_), .A3(new_n723_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n718_), .A2(new_n752_), .B1(new_n751_), .B2(new_n753_), .ZN(G1331gat));
  AOI211_X1 g553(.A(new_n233_), .B(new_n593_), .C1(new_n598_), .C2(new_n600_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n688_), .A2(new_n578_), .A3(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G57gat), .B1(new_n756_), .B2(new_n484_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n655_), .A2(new_n493_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT111), .B1(new_n758_), .B2(new_n233_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n660_), .A2(new_n760_), .A3(new_n234_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n631_), .A2(new_n579_), .A3(new_n640_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n484_), .A2(G57gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n757_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT112), .ZN(G1332gat));
  OAI21_X1  g566(.A(G64gat), .B1(new_n756_), .B2(new_n486_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT48), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n486_), .A2(G64gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n764_), .B2(new_n770_), .ZN(G1333gat));
  NAND4_X1  g570(.A1(new_n688_), .A2(new_n290_), .A3(new_n578_), .A4(new_n755_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(G71gat), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n772_), .B2(G71gat), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n291_), .A2(G71gat), .ZN(new_n777_));
  OAI22_X1  g576(.A1(new_n775_), .A2(new_n776_), .B1(new_n764_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT113), .ZN(G1334gat));
  OAI21_X1  g578(.A(G78gat), .B1(new_n756_), .B2(new_n490_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT50), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n375_), .A2(new_n500_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n764_), .B2(new_n782_), .ZN(G1335gat));
  INV_X1    g582(.A(new_n710_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n579_), .A2(new_n233_), .A3(new_n601_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n634_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G85gat), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n722_), .A2(new_n579_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n484_), .A2(G85gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n788_), .B1(new_n792_), .B2(new_n793_), .ZN(G1336gat));
  NAND2_X1  g593(.A1(new_n786_), .A2(new_n482_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G92gat), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n486_), .A2(G92gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n792_), .B2(new_n797_), .ZN(G1337gat));
  NAND3_X1  g597(.A1(new_n784_), .A2(new_n290_), .A3(new_n785_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G99gat), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n291_), .A2(new_n513_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n791_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n791_), .B2(new_n802_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT51), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n800_), .B(new_n807_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n791_), .A2(new_n518_), .A3(new_n375_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n375_), .B(new_n785_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n518_), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n812_));
  NOR2_X1   g611(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n810_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT53), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n810_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1339gat));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n598_), .A2(new_n600_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n593_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n234_), .A3(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT116), .B1(new_n578_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n755_), .A2(new_n826_), .A3(new_n577_), .A4(new_n576_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n821_), .B1(new_n828_), .B2(new_n632_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT54), .B(new_n631_), .C1(new_n825_), .C2(new_n827_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n233_), .A2(new_n573_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n556_), .A2(new_n559_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(KEYINPUT55), .A3(new_n558_), .A4(new_n547_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n547_), .A2(new_n559_), .A3(new_n556_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n564_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n560_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n560_), .B2(new_n840_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n838_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n833_), .B1(new_n843_), .B2(new_n572_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n560_), .A2(new_n840_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT117), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n560_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n837_), .A4(new_n835_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(KEYINPUT56), .A3(new_n570_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n832_), .B1(new_n844_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n218_), .A2(new_n219_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n219_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n228_), .B1(new_n223_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT118), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n221_), .A2(new_n228_), .A3(new_n224_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n574_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n639_), .B1(new_n850_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT57), .B(new_n639_), .C1(new_n850_), .C2(new_n859_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n857_), .A2(new_n573_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n848_), .A2(KEYINPUT56), .A3(new_n570_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT56), .B1(new_n848_), .B2(new_n570_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(KEYINPUT58), .B(new_n864_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n631_), .A3(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n862_), .A2(new_n863_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n831_), .B1(new_n872_), .B2(new_n640_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n491_), .A2(new_n484_), .A3(new_n291_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n233_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(KEYINPUT59), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n234_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n882_), .B2(new_n877_), .ZN(G1340gat));
  INV_X1    g682(.A(G120gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n579_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n876_), .B(new_n885_), .C1(KEYINPUT60), .C2(new_n884_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n579_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n884_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n876_), .A2(new_n889_), .A3(new_n601_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n640_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1342gat));
  INV_X1    g691(.A(G134gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n876_), .A2(new_n893_), .A3(new_n687_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n632_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n893_), .ZN(G1343gat));
  INV_X1    g695(.A(new_n832_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n687_), .B1(new_n898_), .B2(new_n858_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n870_), .A2(new_n631_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n844_), .A2(new_n849_), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT58), .B1(new_n901_), .B2(new_n864_), .ZN(new_n902_));
  OAI22_X1  g701(.A1(new_n899_), .A2(KEYINPUT57), .B1(new_n900_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n863_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n640_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n831_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n490_), .A2(new_n484_), .A3(new_n482_), .A4(new_n290_), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT119), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910_));
  INV_X1    g709(.A(new_n908_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n873_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n233_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G141gat), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n294_), .B(new_n233_), .C1(new_n909_), .C2(new_n912_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1344gat));
  OAI21_X1  g715(.A(new_n578_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G148gat), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n295_), .B(new_n578_), .C1(new_n909_), .C2(new_n912_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1345gat));
  OAI21_X1  g719(.A(new_n601_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n922_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n601_), .B(new_n924_), .C1(new_n909_), .C2(new_n912_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1346gat));
  NAND2_X1  g725(.A1(new_n705_), .A2(G162gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n907_), .A2(KEYINPUT119), .A3(new_n908_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n910_), .B1(new_n873_), .B2(new_n911_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n687_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n931_));
  INV_X1    g730(.A(G162gat), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1347gat));
  NOR4_X1   g732(.A1(new_n873_), .A2(new_n375_), .A3(new_n486_), .A4(new_n492_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n233_), .A2(new_n252_), .ZN(new_n935_));
  XOR2_X1   g734(.A(new_n935_), .B(KEYINPUT120), .Z(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n492_), .A2(new_n375_), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n907_), .A2(new_n482_), .A3(new_n233_), .A4(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n939_), .A2(new_n940_), .A3(G169gat), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n939_), .B2(G169gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n937_), .B1(new_n941_), .B2(new_n942_), .ZN(G1348gat));
  AOI21_X1  g742(.A(new_n486_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n944_), .A2(new_n578_), .A3(new_n938_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n249_), .A2(KEYINPUT121), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT121), .B(G176gat), .Z(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n945_), .B2(new_n948_), .ZN(G1349gat));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n950_));
  INV_X1    g749(.A(new_n395_), .ZN(new_n951_));
  NAND4_X1  g750(.A1(new_n934_), .A2(new_n950_), .A3(new_n951_), .A4(new_n601_), .ZN(new_n952_));
  AOI21_X1  g751(.A(G183gat), .B1(new_n934_), .B2(new_n601_), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n944_), .A2(new_n951_), .A3(new_n601_), .A4(new_n938_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(KEYINPUT122), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n952_), .B1(new_n953_), .B2(new_n955_), .ZN(G1350gat));
  NAND3_X1  g755(.A1(new_n934_), .A2(new_n396_), .A3(new_n687_), .ZN(new_n957_));
  NAND4_X1  g756(.A1(new_n907_), .A2(new_n482_), .A3(new_n631_), .A4(new_n938_), .ZN(new_n958_));
  AND3_X1   g757(.A1(new_n958_), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n959_));
  AOI21_X1  g758(.A(KEYINPUT123), .B1(new_n958_), .B2(G190gat), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n957_), .B1(new_n959_), .B2(new_n960_), .ZN(G1351gat));
  NOR2_X1   g760(.A1(new_n476_), .A2(new_n290_), .ZN(new_n962_));
  NAND4_X1  g761(.A1(new_n907_), .A2(new_n482_), .A3(new_n233_), .A4(new_n962_), .ZN(new_n963_));
  INV_X1    g762(.A(G197gat), .ZN(new_n964_));
  OAI21_X1  g763(.A(KEYINPUT124), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n963_), .A2(new_n964_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n962_), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n873_), .A2(new_n486_), .A3(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969_));
  NAND4_X1  g768(.A1(new_n968_), .A2(new_n969_), .A3(G197gat), .A4(new_n233_), .ZN(new_n970_));
  AND3_X1   g769(.A1(new_n965_), .A2(new_n966_), .A3(new_n970_), .ZN(G1352gat));
  NAND2_X1  g770(.A1(new_n968_), .A2(new_n578_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g772(.A(new_n640_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n975_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n976_));
  OR3_X1    g775(.A1(new_n975_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977_));
  AOI22_X1  g776(.A1(new_n968_), .A2(new_n974_), .B1(new_n976_), .B2(new_n977_), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n968_), .A2(new_n974_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n979_), .B2(new_n977_), .ZN(G1354gat));
  AND3_X1   g779(.A1(new_n968_), .A2(G218gat), .A3(new_n631_), .ZN(new_n981_));
  NOR4_X1   g780(.A1(new_n873_), .A2(new_n486_), .A3(new_n639_), .A4(new_n967_), .ZN(new_n982_));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983_));
  OR2_X1    g782(.A1(new_n982_), .A2(new_n983_), .ZN(new_n984_));
  AOI21_X1  g783(.A(G218gat), .B1(new_n982_), .B2(new_n983_), .ZN(new_n985_));
  AOI21_X1  g784(.A(new_n981_), .B1(new_n984_), .B2(new_n985_), .ZN(G1355gat));
endmodule


