//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n852_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G204gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(G197gat), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT90), .B1(new_n205_), .B2(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT90), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(new_n203_), .A3(G197gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n204_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n205_), .A2(G204gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT21), .B1(new_n204_), .B2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G211gat), .B(G218gat), .Z(new_n217_));
  AOI21_X1  g016(.A(new_n210_), .B1(new_n217_), .B2(KEYINPUT91), .ZN(new_n218_));
  INV_X1    g017(.A(new_n209_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT91), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT92), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n209_), .B1(new_n220_), .B2(new_n214_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(KEYINPUT92), .A3(new_n218_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n216_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT86), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT3), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n231_), .B(new_n233_), .C1(new_n230_), .C2(new_n228_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT88), .Z(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n232_), .B(KEYINPUT87), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n238_), .B(KEYINPUT1), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n240_), .B(new_n229_), .C1(new_n236_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n227_), .B1(KEYINPUT29), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G78gat), .B(G106gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G228gat), .A2(G233gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(G228gat), .A3(G233gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  OR3_X1    g051(.A1(new_n243_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT28), .B1(new_n243_), .B2(KEYINPUT29), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G22gat), .B(G50gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n253_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .A4(new_n259_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT22), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n268_));
  AOI21_X1  g067(.A(G176gat), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n264_), .B1(new_n269_), .B2(KEYINPUT82), .ZN(new_n270_));
  INV_X1    g069(.A(G176gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n268_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n273_));
  OAI211_X1 g072(.A(KEYINPUT82), .B(new_n271_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT83), .B1(new_n270_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT80), .B(G183gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n277_), .B(KEYINPUT81), .ZN(new_n281_));
  OAI221_X1 g080(.A(new_n279_), .B1(new_n280_), .B2(G190gat), .C1(new_n281_), .C2(new_n278_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT82), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(new_n264_), .A4(new_n274_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n276_), .A2(new_n282_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT84), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT80), .B(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT25), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n290_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n266_), .A2(new_n271_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n296_), .A2(KEYINPUT24), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n277_), .A2(KEYINPUT23), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(new_n281_), .B2(KEYINPUT23), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n296_), .A2(new_n264_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT24), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n295_), .A2(new_n297_), .A3(new_n299_), .A4(new_n301_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n288_), .A2(new_n289_), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n289_), .B1(new_n288_), .B2(new_n302_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT85), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n306_), .B(new_n307_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(KEYINPUT85), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n305_), .B(new_n310_), .Z(new_n311_));
  XOR2_X1   g110(.A(G15gat), .B(G43gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT31), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n311_), .B(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G71gat), .B(G99gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT30), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G227gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  OR2_X1    g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT98), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n243_), .A2(new_n310_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n239_), .A2(new_n309_), .A3(new_n242_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT4), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT4), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n321_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n320_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n324_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT0), .B(G57gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G85gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(G1gat), .B(G29gat), .Z(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n331_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n314_), .A2(new_n318_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n263_), .A2(new_n319_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT27), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT93), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT92), .B1(new_n225_), .B2(new_n218_), .ZN(new_n344_));
  AND4_X1   g143(.A1(KEYINPUT92), .A2(new_n218_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n215_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n303_), .A2(new_n304_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT20), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n343_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT19), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n299_), .B1(G183gat), .B2(G190gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n264_), .B(KEYINPUT95), .Z(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n283_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n279_), .B1(new_n281_), .B2(new_n278_), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(new_n296_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT25), .B(G183gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n290_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n300_), .A2(new_n357_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n355_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n346_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n288_), .A2(new_n302_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT84), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n288_), .A2(new_n289_), .A3(new_n302_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n227_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n349_), .A2(new_n352_), .A3(new_n365_), .A4(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n305_), .A2(new_n227_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT20), .B1(new_n364_), .B2(new_n346_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n351_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G8gat), .B(G36gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT97), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n375_), .A2(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n349_), .A2(new_n351_), .A3(new_n365_), .A4(new_n370_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n352_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n383_), .B1(KEYINPUT100), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n381_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT100), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n342_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n385_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(new_n381_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n393_), .A2(new_n386_), .A3(KEYINPUT27), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n391_), .A2(KEYINPUT101), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT101), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT100), .B1(new_n392_), .B2(new_n381_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n390_), .B1(new_n397_), .B2(new_n388_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT27), .ZN(new_n399_));
  OR3_X1    g198(.A1(new_n393_), .A2(KEYINPUT27), .A3(new_n386_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n396_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n341_), .B1(new_n395_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT102), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT32), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n392_), .B1(new_n404_), .B2(new_n382_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n337_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n382_), .A2(new_n404_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n375_), .A2(KEYINPUT99), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT99), .B1(new_n375_), .B2(new_n407_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n406_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n412_));
  NOR4_X1   g211(.A1(new_n328_), .A2(KEYINPUT33), .A3(new_n330_), .A4(new_n335_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n329_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n324_), .A2(new_n321_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n415_), .A2(new_n336_), .A3(new_n416_), .ZN(new_n417_));
  NOR4_X1   g216(.A1(new_n414_), .A2(new_n393_), .A3(new_n417_), .A4(new_n386_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n263_), .B1(new_n410_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n261_), .A2(new_n262_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n338_), .B(new_n420_), .C1(new_n391_), .C2(new_n394_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n319_), .A2(new_n339_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT101), .B1(new_n391_), .B2(new_n394_), .ZN(new_n425_));
  AOI211_X1 g224(.A(KEYINPUT100), .B(new_n381_), .C1(new_n371_), .C2(new_n374_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n392_), .A2(new_n381_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n389_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n428_), .B2(new_n383_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n396_), .B(new_n400_), .C1(new_n429_), .C2(new_n342_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT102), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n341_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n403_), .A2(new_n424_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G230gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G99gat), .A2(G106gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT66), .ZN(new_n440_));
  OAI22_X1  g239(.A1(new_n440_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  OR4_X1    g240(.A1(new_n440_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G85gat), .B(G92gat), .Z(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT8), .B1(new_n444_), .B2(KEYINPUT67), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(KEYINPUT9), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT9), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(G85gat), .A3(G92gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT10), .B(G99gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT64), .B(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n439_), .A2(new_n448_), .A3(new_n450_), .A4(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n443_), .B(new_n444_), .C1(KEYINPUT67), .C2(KEYINPUT8), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n447_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G57gat), .ZN(new_n457_));
  INV_X1    g256(.A(G64gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G57gat), .A2(G64gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G71gat), .A2(G78gat), .ZN(new_n463_));
  INV_X1    g262(.A(G71gat), .ZN(new_n464_));
  INV_X1    g263(.A(G78gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(new_n463_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT68), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n460_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT68), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n462_), .A2(new_n470_), .A3(new_n463_), .A4(new_n466_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n456_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n456_), .A2(new_n474_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n436_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n477_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT12), .B1(new_n456_), .B2(new_n474_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n483_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n468_), .A2(new_n471_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n469_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT69), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n482_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(KEYINPUT70), .A3(new_n456_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT70), .B1(new_n490_), .B2(new_n456_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n479_), .B(new_n481_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n478_), .B1(new_n494_), .B2(new_n436_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G120gat), .B(G148gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G176gat), .B(G204gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT71), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n495_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(KEYINPUT13), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n504_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G29gat), .B(G36gat), .ZN(new_n508_));
  INV_X1    g307(.A(G43gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(G50gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513_));
  INV_X1    g312(.A(G8gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G8gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  NAND2_X1  g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT76), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n512_), .B(KEYINPUT15), .ZN(new_n521_));
  INV_X1    g320(.A(new_n518_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n520_), .B1(new_n518_), .B2(new_n512_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT77), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n526_), .B1(new_n529_), .B2(new_n525_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(new_n266_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n205_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT79), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n526_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n527_), .B(KEYINPUT77), .ZN(new_n536_));
  INV_X1    g335(.A(new_n525_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT79), .ZN(new_n539_));
  INV_X1    g338(.A(new_n533_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n533_), .B(KEYINPUT78), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n534_), .A2(new_n541_), .B1(new_n530_), .B2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n507_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n434_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT73), .B(G134gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G162gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n512_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n456_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n521_), .A2(new_n456_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  AND2_X1   g359(.A1(new_n560_), .A2(new_n549_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n551_), .B1(new_n561_), .B2(new_n550_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(KEYINPUT74), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n518_), .B(new_n565_), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT75), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n474_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT16), .B(G183gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G211gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(G127gat), .B(G155gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT17), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n566_), .A2(new_n489_), .A3(new_n484_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n566_), .B1(new_n489_), .B2(new_n484_), .ZN(new_n577_));
  OR4_X1    g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .A4(new_n572_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n564_), .A2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n545_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n202_), .B1(new_n582_), .B2(new_n337_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT103), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n562_), .B(new_n563_), .Z(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n564_), .A2(KEYINPUT37), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n579_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n545_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n202_), .A3(new_n337_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT38), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n584_), .A2(new_n594_), .ZN(G1324gat));
  INV_X1    g394(.A(new_n431_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n514_), .B1(new_n582_), .B2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT39), .Z(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n514_), .A3(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(G1325gat));
  INV_X1    g401(.A(G15gat), .ZN(new_n603_));
  INV_X1    g402(.A(new_n423_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n582_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT41), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n592_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1326gat));
  INV_X1    g407(.A(G22gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n582_), .B2(new_n420_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT42), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n592_), .A2(new_n609_), .A3(new_n420_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1327gat));
  AOI21_X1  g412(.A(new_n432_), .B1(new_n431_), .B2(new_n341_), .ZN(new_n614_));
  AOI211_X1 g413(.A(KEYINPUT102), .B(new_n340_), .C1(new_n425_), .C2(new_n430_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n604_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n544_), .A2(new_n580_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n617_), .A2(new_n585_), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(G29gat), .B1(new_n619_), .B2(new_n337_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n564_), .B(new_n586_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT43), .B1(new_n617_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT43), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n587_), .A2(new_n588_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n434_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n618_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT104), .B1(new_n626_), .B2(KEYINPUT44), .ZN(new_n627_));
  INV_X1    g426(.A(new_n618_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n434_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n623_), .B1(new_n434_), .B2(new_n624_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n628_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT44), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n627_), .A2(new_n634_), .B1(KEYINPUT44), .B2(new_n626_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(new_n337_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n620_), .B1(new_n636_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  INV_X1    g437(.A(G36gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n431_), .B(KEYINPUT105), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n619_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT45), .Z(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT44), .B(new_n628_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n626_), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n632_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n596_), .B(new_n644_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n643_), .B1(new_n647_), .B2(G36gat), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n638_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n639_), .B1(new_n635_), .B2(new_n596_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT106), .B(KEYINPUT46), .C1(new_n651_), .C2(new_n643_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n650_), .A2(new_n652_), .ZN(G1329gat));
  NOR2_X1   g452(.A1(new_n423_), .A2(new_n509_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n644_), .B(new_n654_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT107), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n619_), .A2(new_n604_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n509_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n656_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n656_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n655_), .A2(new_n658_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT107), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT47), .B1(new_n665_), .B2(new_n659_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n663_), .A2(new_n666_), .ZN(G1330gat));
  NAND2_X1  g466(.A1(new_n420_), .A2(new_n511_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT109), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n619_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n644_), .A2(new_n420_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n672_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT108), .B1(new_n673_), .B2(G50gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n671_), .B1(new_n627_), .B2(new_n634_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n675_), .A2(new_n676_), .A3(new_n511_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n670_), .B1(new_n674_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT110), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n670_), .C1(new_n674_), .C2(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1331gat));
  INV_X1    g481(.A(new_n507_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n543_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n434_), .A2(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(new_n581_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(G57gat), .A3(new_n337_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n590_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n457_), .B1(new_n689_), .B2(new_n338_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1332gat));
  AOI21_X1  g490(.A(new_n458_), .B1(new_n687_), .B2(new_n641_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT48), .Z(new_n693_));
  NOR2_X1   g492(.A1(new_n640_), .A2(G64gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT111), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n689_), .B2(new_n695_), .ZN(G1333gat));
  AOI21_X1  g495(.A(new_n464_), .B1(new_n687_), .B2(new_n604_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT49), .Z(new_n698_));
  NOR2_X1   g497(.A1(new_n423_), .A2(G71gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT112), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n689_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT113), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(G1334gat));
  AOI21_X1  g502(.A(new_n465_), .B1(new_n687_), .B2(new_n420_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT50), .Z(new_n705_));
  NAND2_X1  g504(.A1(new_n420_), .A2(new_n465_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n689_), .B2(new_n706_), .ZN(G1335gat));
  NAND2_X1  g506(.A1(new_n685_), .A2(new_n580_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n617_), .A2(new_n585_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n337_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n337_), .A2(G85gat), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT114), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n711_), .B2(new_n713_), .ZN(G1336gat));
  AOI21_X1  g513(.A(G92gat), .B1(new_n709_), .B2(new_n596_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n711_), .A2(new_n641_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(G92gat), .ZN(G1337gat));
  NAND2_X1  g516(.A1(new_n711_), .A2(new_n604_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n604_), .A2(new_n451_), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n718_), .A2(G99gat), .B1(new_n709_), .B2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT51), .Z(G1338gat));
  NAND2_X1  g520(.A1(new_n711_), .A2(new_n420_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(G106gat), .A3(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n709_), .A2(new_n452_), .A3(new_n420_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n725_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n726_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n494_), .B2(new_n436_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT116), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n490_), .A2(new_n456_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT70), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  AOI211_X1 g535(.A(new_n477_), .B(new_n480_), .C1(new_n736_), .C2(new_n491_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n733_), .B1(new_n737_), .B2(new_n435_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n494_), .A2(KEYINPUT116), .A3(new_n436_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n732_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT55), .B1(new_n737_), .B2(new_n435_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT116), .B1(new_n494_), .B2(new_n436_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n737_), .A2(new_n733_), .A3(new_n435_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n500_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT56), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n740_), .A2(new_n744_), .A3(KEYINPUT56), .A4(new_n500_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n495_), .A2(new_n500_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(new_n684_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n524_), .A2(new_n537_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n540_), .B1(new_n536_), .B2(new_n525_), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n534_), .A2(new_n541_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n503_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n564_), .B1(new_n752_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(KEYINPUT117), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT117), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT57), .B1(new_n757_), .B2(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT119), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n745_), .A2(new_n764_), .A3(new_n746_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n748_), .B(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n755_), .B(new_n751_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT120), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT58), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT58), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(KEYINPUT120), .A3(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n624_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n579_), .B1(new_n763_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n589_), .A2(new_n507_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n543_), .ZN(new_n779_));
  NOR4_X1   g578(.A1(new_n589_), .A2(KEYINPUT54), .A3(new_n507_), .A4(new_n684_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n337_), .B(new_n263_), .C1(new_n776_), .C2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n596_), .A2(new_n423_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G113gat), .B1(new_n785_), .B2(new_n684_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT59), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n778_), .A2(new_n543_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT54), .ZN(new_n790_));
  INV_X1    g589(.A(new_n780_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n770_), .A2(KEYINPUT120), .A3(new_n773_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n773_), .B1(new_n770_), .B2(KEYINPUT120), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n621_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n760_), .A2(new_n762_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n580_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n420_), .B1(new_n792_), .B2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n798_), .A2(KEYINPUT59), .A3(new_n337_), .A4(new_n783_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n788_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n684_), .A2(G113gat), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT121), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n786_), .B1(new_n800_), .B2(new_n802_), .ZN(G1340gat));
  INV_X1    g602(.A(G120gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n683_), .B2(KEYINPUT60), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n785_), .B(new_n805_), .C1(KEYINPUT60), .C2(new_n804_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n683_), .B1(new_n788_), .B2(new_n799_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n804_), .ZN(G1341gat));
  AOI21_X1  g607(.A(G127gat), .B1(new_n785_), .B2(new_n579_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n800_), .A2(G127gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n579_), .ZN(G1342gat));
  XOR2_X1   g610(.A(KEYINPUT122), .B(G134gat), .Z(new_n812_));
  NOR2_X1   g611(.A1(new_n621_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n800_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n785_), .A2(new_n564_), .ZN(new_n816_));
  INV_X1    g615(.A(G134gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(new_n815_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n813_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n788_), .B2(new_n799_), .ZN(new_n821_));
  AOI21_X1  g620(.A(G134gat), .B1(new_n785_), .B2(new_n564_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT123), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(new_n823_), .ZN(G1343gat));
  AOI21_X1  g623(.A(new_n641_), .B1(new_n792_), .B2(new_n797_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n604_), .A2(new_n263_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n338_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n684_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n507_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g633(.A1(new_n829_), .A2(new_n580_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT61), .B(G155gat), .Z(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1346gat));
  AOI21_X1  g636(.A(G162gat), .B1(new_n830_), .B2(new_n564_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n829_), .A2(new_n621_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(G162gat), .B2(new_n839_), .ZN(G1347gat));
  NAND2_X1  g639(.A1(new_n792_), .A2(new_n797_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(new_n341_), .A3(new_n641_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G169gat), .B1(new_n842_), .B2(new_n543_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n842_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(new_n684_), .C1(new_n273_), .C2(new_n272_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n844_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n847_), .A3(new_n848_), .ZN(G1348gat));
  NOR2_X1   g648(.A1(new_n842_), .A2(new_n683_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n271_), .ZN(G1349gat));
  NOR2_X1   g650(.A1(new_n842_), .A2(new_n580_), .ZN(new_n852_));
  MUX2_X1   g651(.A(new_n280_), .B(new_n360_), .S(new_n852_), .Z(G1350gat));
  NAND3_X1  g652(.A1(new_n846_), .A2(new_n564_), .A3(new_n290_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G190gat), .B1(new_n842_), .B2(new_n621_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(KEYINPUT124), .A3(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1351gat));
  XNOR2_X1  g659(.A(KEYINPUT126), .B(G197gat), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n827_), .A2(new_n337_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n641_), .B(new_n865_), .C1(new_n776_), .C2(new_n781_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n863_), .A2(new_n864_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n861_), .B1(new_n869_), .B2(new_n543_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n868_), .A2(KEYINPUT126), .A3(new_n205_), .A4(new_n684_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1352gat));
  NAND2_X1  g671(.A1(new_n868_), .A2(new_n507_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g673(.A1(new_n868_), .A2(new_n579_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n876_));
  AND2_X1   g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n875_), .B2(new_n876_), .ZN(G1354gat));
  INV_X1    g678(.A(G218gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n868_), .B2(new_n624_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT127), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n866_), .A2(G218gat), .A3(new_n585_), .A4(new_n867_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(new_n883_), .A3(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT127), .B1(new_n881_), .B2(new_n884_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1355gat));
endmodule


