//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT72), .B(G15gat), .ZN(new_n206_));
  INV_X1    g005(.A(G22gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G1gat), .B(G8gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n212_), .B(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n205_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n204_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT79), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n212_), .B(new_n213_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n204_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  AND4_X1   g025(.A1(KEYINPUT78), .A2(new_n226_), .A3(G229gat), .A4(G233gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n219_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT78), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n221_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G141gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G169gat), .B(G197gat), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n231_), .B(new_n232_), .Z(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n221_), .B(new_n233_), .C1(new_n227_), .C2(new_n229_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G226gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT19), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT20), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G183gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(KEYINPUT23), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n245_), .A2(G190gat), .B1(KEYINPUT23), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G169gat), .ZN(new_n248_));
  INV_X1    g047(.A(G176gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(KEYINPUT24), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT95), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(KEYINPUT23), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT23), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(G183gat), .A3(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT95), .ZN(new_n257_));
  OR3_X1    g056(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT25), .B(G183gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G190gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n260_), .A2(new_n261_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n252_), .A2(new_n259_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n248_), .A2(KEYINPUT22), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(G169gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT96), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n249_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n264_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n255_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n254_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n276_), .A2(new_n277_), .B1(KEYINPUT23), .B2(new_n246_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n266_), .B1(new_n274_), .B2(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(G197gat), .A2(G204gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G197gat), .A2(G204gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(KEYINPUT21), .A3(new_n283_), .ZN(new_n287_));
  INV_X1    g086(.A(G218gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G211gat), .ZN(new_n289_));
  INV_X1    g088(.A(G211gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G218gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT92), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n289_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n292_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n286_), .B(new_n287_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n295_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n287_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(new_n293_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n243_), .B1(new_n281_), .B2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n296_), .A2(new_n299_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n244_), .A2(KEYINPUT25), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G183gat), .ZN(new_n305_));
  INV_X1    g104(.A(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT26), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G190gat), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n303_), .A2(new_n305_), .A3(new_n307_), .A4(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT80), .ZN(new_n311_));
  AND2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n262_), .B2(new_n312_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n250_), .A2(KEYINPUT80), .A3(KEYINPUT24), .A4(new_n264_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT81), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n310_), .A2(new_n313_), .A3(new_n314_), .A4(KEYINPUT81), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n276_), .A2(new_n277_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n253_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n317_), .A2(new_n318_), .A3(new_n320_), .A4(new_n258_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n279_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n322_), .A2(KEYINPUT83), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(KEYINPUT83), .ZN(new_n324_));
  NOR2_X1   g123(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G169gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n323_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n302_), .B1(new_n321_), .B2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n301_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n320_), .B1(G183gat), .B2(G190gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n268_), .A2(G169gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n248_), .A2(KEYINPUT22), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT96), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n312_), .B1(new_n335_), .B2(new_n249_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n257_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n250_), .A2(KEYINPUT24), .A3(new_n264_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n310_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n330_), .A2(new_n336_), .B1(new_n340_), .B2(new_n259_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT97), .B1(new_n341_), .B2(new_n302_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n321_), .A2(new_n302_), .A3(new_n327_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT97), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n281_), .A2(new_n344_), .A3(new_n300_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n342_), .A2(KEYINPUT20), .A3(new_n343_), .A4(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n241_), .B(KEYINPUT94), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n329_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  AOI211_X1 g153(.A(new_n352_), .B(new_n329_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n239_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n346_), .A2(new_n347_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n329_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n353_), .A3(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n273_), .B(new_n264_), .C1(new_n279_), .C2(new_n278_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n360_), .A2(KEYINPUT102), .A3(new_n266_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT102), .B1(new_n360_), .B2(new_n266_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n361_), .A2(new_n362_), .A3(new_n300_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n324_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n326_), .B1(new_n322_), .B2(KEYINPUT83), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n318_), .A2(new_n320_), .A3(new_n258_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n317_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n365_), .B1(new_n370_), .B2(new_n302_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n241_), .B1(new_n363_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n281_), .A2(new_n300_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n242_), .B1(new_n373_), .B2(KEYINPUT97), .ZN(new_n374_));
  INV_X1    g173(.A(new_n347_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n343_), .A4(new_n345_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n353_), .B1(new_n372_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT103), .ZN(new_n378_));
  OAI211_X1 g177(.A(KEYINPUT27), .B(new_n359_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  AOI211_X1 g178(.A(KEYINPUT103), .B(new_n353_), .C1(new_n372_), .C2(new_n376_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n356_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(G78gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G106gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  OR3_X1    g187(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n389_), .A2(new_n390_), .B1(G155gat), .B2(G162gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT88), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n394_), .A2(G141gat), .A3(G148gat), .ZN(new_n395_));
  INV_X1    g194(.A(G141gat), .ZN(new_n396_));
  INV_X1    g195(.A(G148gat), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n393_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n392_), .B2(KEYINPUT88), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n391_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT3), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n394_), .B1(G141gat), .B2(G148gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G141gat), .A2(G148gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT2), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n407_), .A2(new_n412_), .A3(new_n400_), .A4(new_n393_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(KEYINPUT89), .A3(new_n391_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n404_), .A2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G141gat), .B(G148gat), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n389_), .A2(new_n390_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  OR3_X1    g217(.A1(new_n418_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT87), .B1(new_n418_), .B2(KEYINPUT1), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(KEYINPUT1), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT86), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n416_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n388_), .B1(new_n415_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n387_), .B1(new_n426_), .B2(new_n302_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n422_), .B(KEYINPUT86), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n428_), .A2(new_n417_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n404_), .A2(new_n414_), .B1(new_n429_), .B2(new_n416_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n300_), .B(new_n386_), .C1(new_n430_), .C2(new_n388_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(KEYINPUT91), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT93), .ZN(new_n433_));
  XOR2_X1   g232(.A(G22gat), .B(G50gat), .Z(new_n434_));
  AND3_X1   g233(.A1(new_n413_), .A2(KEYINPUT89), .A3(new_n391_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT89), .B1(new_n413_), .B2(new_n391_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n425_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n434_), .B1(new_n437_), .B2(KEYINPUT29), .ZN(new_n438_));
  INV_X1    g237(.A(new_n434_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n430_), .A2(new_n388_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n438_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT93), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n427_), .A2(new_n447_), .A3(new_n431_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n433_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n432_), .A2(new_n443_), .A3(KEYINPUT93), .A4(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n382_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n453_), .B(G15gat), .Z(new_n454_));
  XOR2_X1   g253(.A(new_n454_), .B(KEYINPUT30), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n370_), .B(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G127gat), .B(G134gat), .Z(new_n457_));
  XOR2_X1   g256(.A(G113gat), .B(G120gat), .Z(new_n458_));
  XOR2_X1   g257(.A(new_n457_), .B(new_n458_), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT31), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT84), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n461_), .B2(new_n460_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n456_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G71gat), .B(G99gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G43gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n466_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n437_), .A2(new_n459_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n415_), .A2(new_n460_), .A3(new_n425_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT4), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT4), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n437_), .A2(new_n473_), .A3(new_n459_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G225gat), .A2(G233gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G1gat), .B(G29gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(G57gat), .B(G85gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n477_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n478_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n476_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n483_), .B1(new_n488_), .B2(new_n485_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n469_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n452_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n372_), .A2(new_n376_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT32), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n352_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT100), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n494_), .A2(new_n496_), .B1(new_n348_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n490_), .A2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT33), .B(new_n483_), .C1(new_n488_), .C2(new_n485_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT99), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT33), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n489_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n357_), .A2(new_n358_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n352_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n470_), .A2(new_n471_), .A3(new_n477_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n484_), .B(new_n506_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n503_), .A2(new_n359_), .A3(new_n505_), .A4(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n499_), .B1(new_n501_), .B2(new_n508_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n360_), .A2(new_n266_), .B1(new_n299_), .B2(new_n296_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT20), .B1(new_n510_), .B2(new_n344_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n281_), .A2(new_n344_), .A3(new_n300_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n321_), .A2(new_n302_), .A3(new_n327_), .ZN(new_n513_));
  NOR4_X1   g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .A4(new_n347_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n241_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n328_), .A2(new_n364_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT102), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n281_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n360_), .A2(KEYINPUT102), .A3(new_n266_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n302_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n515_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n352_), .B1(new_n514_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT103), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n377_), .A2(new_n378_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n239_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n449_), .A2(new_n450_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n356_), .A4(new_n491_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n509_), .A2(new_n451_), .B1(new_n528_), .B2(KEYINPUT104), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n449_), .A2(new_n487_), .A3(new_n489_), .A4(new_n450_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT104), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n356_), .A4(new_n526_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n469_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n493_), .B1(new_n534_), .B2(KEYINPUT105), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT104), .B1(new_n381_), .B2(new_n530_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n490_), .A2(new_n498_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n505_), .A2(new_n359_), .A3(new_n507_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n489_), .A2(new_n502_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT99), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n500_), .B(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n537_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n536_), .B(new_n533_), .C1(new_n543_), .C2(new_n527_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n469_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT105), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n238_), .B1(new_n535_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550_));
  XOR2_X1   g349(.A(G85gat), .B(G92gat), .Z(new_n551_));
  NOR2_X1   g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT6), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n551_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT8), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n557_), .B1(KEYINPUT9), .B2(new_n551_), .ZN(new_n561_));
  XOR2_X1   g360(.A(KEYINPUT10), .B(G99gat), .Z(new_n562_));
  INV_X1    g361(.A(G106gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT65), .B(G85gat), .ZN(new_n565_));
  INV_X1    g364(.A(G92gat), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n565_), .A2(KEYINPUT9), .A3(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n561_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n560_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n217_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT34), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n558_), .B(KEYINPUT8), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT67), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT67), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n560_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n568_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  OAI221_X1 g376(.A(new_n570_), .B1(KEYINPUT35), .B2(new_n572_), .C1(new_n577_), .C2(new_n205_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n570_), .ZN(new_n580_));
  OAI211_X1 g379(.A(KEYINPUT35), .B(new_n572_), .C1(new_n580_), .C2(KEYINPUT69), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n581_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT70), .ZN(new_n586_));
  XOR2_X1   g385(.A(G134gat), .B(G162gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT36), .Z(new_n589_));
  AND2_X1   g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n582_), .A2(new_n591_), .A3(new_n583_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n549_), .B(new_n550_), .C1(new_n590_), .C2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n584_), .A2(new_n589_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(KEYINPUT71), .A2(KEYINPUT37), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n549_), .A2(new_n550_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n595_), .A2(new_n592_), .A3(new_n596_), .A4(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT64), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n604_));
  XOR2_X1   g403(.A(G71gat), .B(G78gat), .Z(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n569_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT66), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n569_), .A2(KEYINPUT66), .A3(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n569_), .A2(new_n609_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n602_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n569_), .B2(new_n609_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n602_), .B1(new_n569_), .B2(new_n609_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n609_), .A2(new_n617_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n618_), .B(new_n619_), .C1(new_n577_), .C2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G120gat), .B(G148gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT5), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n622_), .B(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT13), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(KEYINPUT68), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n628_), .A2(KEYINPUT68), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n631_), .B2(new_n629_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n609_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT73), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(new_n222_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G127gat), .B(G155gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT17), .Z(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT75), .B1(new_n637_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(KEYINPUT17), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(new_n637_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n637_), .A2(KEYINPUT75), .A3(new_n643_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(KEYINPUT76), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT76), .B1(new_n646_), .B2(new_n647_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n600_), .A2(new_n633_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n548_), .A2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(G1gat), .A3(new_n491_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n590_), .A2(new_n593_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n535_), .B2(new_n547_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n633_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n646_), .A2(new_n647_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n659_), .A2(new_n238_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n658_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n491_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n654_), .A2(new_n655_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n656_), .A2(new_n664_), .A3(new_n665_), .ZN(G1324gat));
  OAI21_X1  g465(.A(G8gat), .B1(new_n663_), .B2(new_n382_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT39), .ZN(new_n668_));
  INV_X1    g467(.A(new_n653_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n210_), .A3(new_n381_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT40), .Z(G1325gat));
  NOR3_X1   g471(.A1(new_n653_), .A2(G15gat), .A3(new_n545_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT107), .ZN(new_n674_));
  OAI21_X1  g473(.A(G15gat), .B1(new_n663_), .B2(new_n545_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT41), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(KEYINPUT41), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n676_), .A3(new_n677_), .ZN(G1326gat));
  OR2_X1    g477(.A1(new_n451_), .A2(KEYINPUT108), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n451_), .A2(KEYINPUT108), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G22gat), .B1(new_n663_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT42), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n669_), .A2(new_n207_), .A3(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(new_n650_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n657_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(new_n659_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n548_), .A2(new_n689_), .ZN(new_n690_));
  OR3_X1    g489(.A1(new_n690_), .A2(G29gat), .A3(new_n491_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n544_), .A2(KEYINPUT105), .A3(new_n545_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n493_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n692_), .B(new_n599_), .C1(new_n695_), .C2(new_n546_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n600_), .B1(new_n535_), .B2(new_n547_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n659_), .A2(new_n650_), .A3(new_n238_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(KEYINPUT44), .A3(new_n701_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n490_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT110), .ZN(new_n708_));
  OAI21_X1  g507(.A(G29gat), .B1(new_n707_), .B2(KEYINPUT110), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n691_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  NOR3_X1   g509(.A1(new_n690_), .A2(G36gat), .A3(new_n382_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT45), .Z(new_n712_));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n704_), .A2(new_n381_), .A3(new_n705_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n712_), .B(KEYINPUT46), .C1(new_n714_), .C2(new_n713_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1329gat));
  NAND3_X1  g518(.A1(new_n706_), .A2(G43gat), .A3(new_n469_), .ZN(new_n720_));
  INV_X1    g519(.A(G43gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n690_), .B2(new_n545_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n720_), .A2(KEYINPUT47), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT47), .B1(new_n720_), .B2(new_n722_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1330gat));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n706_), .A2(new_n527_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G50gat), .ZN(new_n728_));
  INV_X1    g527(.A(G50gat), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT111), .B(new_n729_), .C1(new_n706_), .C2(new_n527_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n681_), .A2(new_n729_), .ZN(new_n731_));
  OAI22_X1  g530(.A1(new_n728_), .A2(new_n730_), .B1(new_n690_), .B2(new_n731_), .ZN(G1331gat));
  AOI21_X1  g531(.A(new_n237_), .B1(new_n535_), .B2(new_n547_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n687_), .A2(new_n599_), .A3(new_n633_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT112), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n491_), .B1(new_n735_), .B2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G57gat), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n687_), .A2(new_n237_), .A3(new_n633_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n658_), .A2(G57gat), .A3(new_n490_), .A4(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT113), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n740_), .A2(new_n743_), .ZN(G1332gat));
  NAND2_X1  g543(.A1(new_n658_), .A2(new_n741_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G64gat), .B1(new_n745_), .B2(new_n382_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT48), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n735_), .A2(G64gat), .A3(new_n382_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT114), .Z(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n745_), .B2(new_n545_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n545_), .A2(G71gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n735_), .B2(new_n753_), .ZN(G1334gat));
  OAI21_X1  g553(.A(G78gat), .B1(new_n745_), .B2(new_n682_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n736_), .A2(new_n384_), .A3(new_n681_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1335gat));
  NAND4_X1  g557(.A1(new_n733_), .A2(new_n659_), .A3(new_n687_), .A4(new_n657_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n490_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n650_), .A2(new_n633_), .A3(new_n237_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n599_), .B1(new_n695_), .B2(new_n546_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n698_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n765_), .B2(new_n696_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n491_), .A2(new_n565_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n761_), .B1(new_n766_), .B2(new_n767_), .ZN(G1336gat));
  NAND2_X1  g567(.A1(new_n700_), .A2(new_n762_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G92gat), .B1(new_n769_), .B2(new_n382_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n760_), .A2(new_n566_), .A3(new_n381_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n769_), .B2(new_n545_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n760_), .A2(new_n469_), .A3(new_n562_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n775_), .B(new_n776_), .Z(G1338gat));
  NAND3_X1  g576(.A1(new_n760_), .A2(new_n563_), .A3(new_n527_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n451_), .B(new_n763_), .C1(new_n765_), .C2(new_n696_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n563_), .B1(new_n780_), .B2(KEYINPUT116), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n769_), .B2(new_n451_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n779_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n700_), .A2(KEYINPUT116), .A3(new_n527_), .A4(new_n762_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT116), .B1(new_n766_), .B2(new_n527_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(KEYINPUT52), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n778_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n778_), .C1(new_n784_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  XNOR2_X1  g592(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n651_), .B2(new_n237_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n687_), .A2(new_n599_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n797_), .A2(new_n238_), .A3(new_n633_), .A4(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n622_), .A2(new_n626_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n618_), .B1(new_n577_), .B2(new_n620_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n602_), .B1(new_n614_), .B2(new_n803_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n577_), .A2(new_n620_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n805_), .A2(KEYINPUT55), .A3(new_n618_), .A4(new_n619_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n621_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n804_), .A2(new_n806_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n626_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT118), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n809_), .A2(new_n814_), .A3(new_n626_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .A4(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n809_), .A2(KEYINPUT56), .A3(new_n626_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n810_), .B2(KEYINPUT118), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n812_), .B1(new_n819_), .B2(new_n815_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n802_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n226_), .A2(new_n220_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n220_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n233_), .B1(new_n216_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT120), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n826_), .A2(new_n236_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n627_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n821_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n800_), .B1(new_n829_), .B2(new_n657_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n657_), .B1(new_n821_), .B2(new_n828_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT57), .ZN(new_n832_));
  INV_X1    g631(.A(new_n801_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n810_), .A2(new_n813_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n817_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n827_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n827_), .A2(KEYINPUT58), .A3(new_n833_), .A4(new_n835_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n599_), .A3(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n830_), .A2(new_n832_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n799_), .B1(new_n841_), .B2(new_n661_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n452_), .A2(new_n545_), .A3(new_n491_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT59), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n840_), .B1(new_n831_), .B2(KEYINPUT57), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n831_), .A2(KEYINPUT57), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n687_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n796_), .A2(new_n798_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(new_n843_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n845_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n237_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G113gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n842_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n843_), .ZN(new_n857_));
  OR3_X1    g656(.A1(new_n857_), .A2(G113gat), .A3(new_n238_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(G1340gat));
  XOR2_X1   g658(.A(KEYINPUT121), .B(G120gat), .Z(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n633_), .B2(KEYINPUT60), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT122), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n863_));
  INV_X1    g662(.A(new_n860_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n856_), .A2(new_n843_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n853_), .B2(new_n659_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n845_), .A2(new_n852_), .A3(new_n869_), .A4(new_n659_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n864_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n870_), .B2(new_n872_), .ZN(G1341gat));
  NAND2_X1  g672(.A1(new_n853_), .A2(new_n660_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G127gat), .ZN(new_n875_));
  OR3_X1    g674(.A1(new_n857_), .A2(G127gat), .A3(new_n687_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1342gat));
  NAND2_X1  g676(.A1(new_n853_), .A2(new_n599_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G134gat), .ZN(new_n879_));
  OR4_X1    g678(.A1(G134gat), .A2(new_n857_), .A3(new_n593_), .A4(new_n590_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1343gat));
  NOR2_X1   g680(.A1(new_n842_), .A2(new_n469_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n381_), .A2(new_n491_), .A3(new_n451_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n238_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n396_), .ZN(G1344gat));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n633_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n397_), .ZN(G1345gat));
  NOR2_X1   g687(.A1(new_n884_), .A2(new_n687_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT61), .B(G155gat), .Z(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1346gat));
  INV_X1    g690(.A(G162gat), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n884_), .A2(new_n892_), .A3(new_n600_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n882_), .A2(new_n657_), .A3(new_n883_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n892_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT125), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n897_), .A3(new_n892_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n893_), .B1(new_n896_), .B2(new_n898_), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n492_), .A2(new_n382_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n681_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n850_), .A2(new_n335_), .A3(new_n237_), .A4(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n902_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n238_), .B(new_n904_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n903_), .B(KEYINPUT62), .C1(new_n905_), .C2(new_n248_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n850_), .A2(new_n902_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n907_), .B(G169gat), .C1(new_n908_), .C2(new_n238_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT126), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n906_), .A2(new_n912_), .A3(new_n909_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1348gat));
  INV_X1    g713(.A(new_n908_), .ZN(new_n915_));
  AOI21_X1  g714(.A(G176gat), .B1(new_n915_), .B2(new_n659_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n842_), .A2(new_n527_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n633_), .A2(new_n249_), .A3(new_n901_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(G1349gat));
  NOR3_X1   g718(.A1(new_n908_), .A2(new_n260_), .A3(new_n661_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(new_n650_), .A3(new_n900_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n244_), .B2(new_n921_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n908_), .B2(new_n600_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n657_), .A2(new_n261_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n908_), .B2(new_n924_), .ZN(G1351gat));
  NOR2_X1   g724(.A1(new_n382_), .A2(new_n530_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n882_), .A2(new_n237_), .A3(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g727(.A1(new_n882_), .A2(new_n926_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n633_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n931_), .A2(G204gat), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(G204gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n930_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(new_n930_), .B2(new_n933_), .ZN(G1353gat));
  INV_X1    g734(.A(new_n929_), .ZN(new_n936_));
  XOR2_X1   g735(.A(KEYINPUT63), .B(G211gat), .Z(new_n937_));
  NAND3_X1  g736(.A1(new_n936_), .A2(new_n660_), .A3(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n939_), .B1(new_n929_), .B2(new_n661_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1354gat));
  OAI21_X1  g740(.A(G218gat), .B1(new_n929_), .B2(new_n600_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n657_), .A2(new_n288_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n929_), .B2(new_n943_), .ZN(G1355gat));
endmodule


