//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n596_, new_n597_, new_n598_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT3), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT2), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT85), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT83), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n211_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT84), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n217_), .B(new_n214_), .C1(KEYINPUT1), .C2(new_n212_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n206_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n208_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n205_), .B1(new_n215_), .B2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n211_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n220_), .A3(new_n204_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(KEYINPUT4), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G225gat), .A2(G233gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT93), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n205_), .B(new_n229_), .C1(new_n215_), .C2(new_n221_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n222_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G1gat), .B(G29gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(G85gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT0), .B(G57gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n232_), .A2(KEYINPUT96), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT96), .B1(new_n232_), .B2(new_n237_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n231_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT97), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(KEYINPUT97), .B(new_n231_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G226gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT19), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G197gat), .B(G204gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT21), .B(new_n247_), .C1(new_n249_), .C2(KEYINPUT87), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n250_), .B(new_n251_), .C1(KEYINPUT21), .C2(new_n249_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT21), .A3(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT23), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(G183gat), .B2(G190gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT90), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT22), .B(G169gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT89), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n260_), .B(new_n261_), .C1(G176gat), .C2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT25), .B(G183gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G190gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G169gat), .ZN(new_n268_));
  INV_X1    g067(.A(G176gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT24), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(KEYINPUT24), .A3(new_n261_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n267_), .A2(new_n258_), .A3(new_n271_), .A4(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n256_), .B1(new_n264_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G169gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n259_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n273_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n255_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT20), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n245_), .B1(new_n277_), .B2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G8gat), .B(G36gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  AOI21_X1  g090(.A(new_n283_), .B1(new_n255_), .B2(new_n281_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n264_), .A2(new_n273_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n292_), .B1(new_n293_), .B2(new_n255_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(new_n245_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n286_), .A2(new_n291_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n291_), .B1(new_n286_), .B2(new_n296_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n242_), .A2(new_n243_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT95), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n222_), .A2(KEYINPUT4), .A3(new_n224_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n230_), .A2(new_n227_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n222_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n225_), .A2(KEYINPUT95), .A3(new_n227_), .A4(new_n230_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n305_), .A2(new_n236_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT33), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n237_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n308_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n293_), .A2(new_n255_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT91), .ZN(new_n316_));
  INV_X1    g115(.A(new_n245_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n276_), .A4(new_n284_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n294_), .A2(new_n245_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n286_), .A2(new_n296_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n291_), .A2(KEYINPUT32), .ZN(new_n322_));
  MUX2_X1   g121(.A(new_n320_), .B(new_n321_), .S(new_n322_), .Z(new_n323_));
  OAI22_X1  g122(.A1(new_n301_), .A2(new_n310_), .B1(new_n314_), .B2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n215_), .A2(new_n221_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n255_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT86), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G228gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n328_), .A2(G228gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(G233gat), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n255_), .B(new_n332_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G78gat), .B(G106gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT88), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n325_), .A2(new_n326_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT28), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n341_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n334_), .A2(new_n335_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n336_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n338_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n348_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n324_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT27), .B1(new_n298_), .B2(new_n300_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n286_), .A2(new_n296_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n291_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n355_), .A2(KEYINPUT99), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT98), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n320_), .B2(new_n356_), .ZN(new_n359_));
  AOI211_X1 g158(.A(KEYINPUT98), .B(new_n291_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n357_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT27), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n298_), .B2(KEYINPUT99), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n354_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n313_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n353_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(G15gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G43gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n373_), .A2(KEYINPUT81), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(KEYINPUT81), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n281_), .B(KEYINPUT30), .Z(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n377_), .B(new_n378_), .C1(new_n374_), .C2(new_n376_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n379_), .A2(KEYINPUT31), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(KEYINPUT31), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n204_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n205_), .A3(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n361_), .A2(new_n363_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n354_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(new_n351_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n385_), .A2(new_n313_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n367_), .A2(new_n385_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G85gat), .A2(G92gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT9), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G85gat), .A2(G92gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT65), .B1(new_n398_), .B2(new_n395_), .ZN(new_n399_));
  AND2_X1   g198(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n400_));
  NOR2_X1   g199(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT65), .B(new_n395_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n397_), .B1(new_n399_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT66), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n395_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT65), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n396_), .B1(new_n408_), .B2(new_n402_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT10), .B(G99gat), .Z(new_n412_));
  INV_X1    g211(.A(G106gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G99gat), .A2(G106gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT6), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(G99gat), .A3(G106gat), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n412_), .A2(new_n413_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n405_), .A2(new_n411_), .A3(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G29gat), .B(G36gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G43gat), .B(G50gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT8), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT68), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n416_), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n414_), .A2(KEYINPUT6), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n415_), .A2(new_n417_), .A3(KEYINPUT68), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT69), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G99gat), .A2(G106gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n432_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n430_), .B(new_n433_), .C1(new_n436_), .C2(new_n431_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT67), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n431_), .B1(new_n440_), .B2(new_n432_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n431_), .A2(new_n432_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT69), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n429_), .A2(new_n437_), .A3(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n393_), .A2(new_n395_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n423_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n423_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n441_), .A2(new_n442_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n415_), .A2(new_n417_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n419_), .B(new_n422_), .C1(new_n446_), .C2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G232gat), .A2(G233gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT34), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT35), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n451_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n404_), .A2(KEYINPUT66), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n418_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n459_));
  OAI22_X1  g258(.A1(new_n446_), .A2(new_n450_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n422_), .B(KEYINPUT15), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n460_), .A2(KEYINPUT72), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT72), .B1(new_n460_), .B2(new_n461_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n457_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n454_), .A2(new_n455_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  OAI221_X1 g265(.A(new_n457_), .B1(new_n455_), .B2(new_n454_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G190gat), .B(G218gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G134gat), .B(G162gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT74), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n466_), .A2(new_n467_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT75), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT75), .A4(new_n473_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n466_), .A2(new_n467_), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n470_), .B(KEYINPUT36), .Z(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(KEYINPUT76), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT37), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT77), .B(G1gat), .Z(new_n485_));
  INV_X1    g284(.A(G8gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G8gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G231gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT78), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n494_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n499_));
  XOR2_X1   g298(.A(G71gat), .B(G78gat), .Z(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n499_), .A2(new_n500_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n501_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n497_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G127gat), .B(G155gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT16), .ZN(new_n510_));
  XOR2_X1   g309(.A(G183gat), .B(G211gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n507_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n508_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n506_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n476_), .A2(new_n477_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT76), .A3(KEYINPUT37), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n484_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT13), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT71), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n520_), .A2(KEYINPUT71), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G120gat), .B(G148gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT5), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G176gat), .B(G204gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n505_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n419_), .B(new_n527_), .C1(new_n446_), .C2(new_n450_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G230gat), .A2(G233gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n444_), .A2(new_n445_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n450_), .B1(new_n531_), .B2(KEYINPUT8), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n458_), .A2(new_n459_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n505_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT12), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n460_), .A2(new_n536_), .A3(new_n505_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n530_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n529_), .B1(new_n534_), .B2(new_n528_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n526_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n528_), .A2(new_n529_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n460_), .A2(new_n536_), .A3(new_n505_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n536_), .B1(new_n460_), .B2(new_n505_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n539_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n526_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n540_), .A2(KEYINPUT70), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT70), .B1(new_n540_), .B2(new_n547_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n521_), .B(new_n522_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT70), .ZN(new_n551_));
  INV_X1    g350(.A(new_n547_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n546_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n540_), .A2(KEYINPUT70), .A3(new_n547_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n554_), .A2(KEYINPUT71), .A3(new_n520_), .A4(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n519_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n558_), .A2(KEYINPUT79), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(KEYINPUT79), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n494_), .B(new_n422_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n461_), .A2(new_n493_), .A3(new_n492_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n494_), .B2(new_n422_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n561_), .A2(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G169gat), .B(G197gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  OR2_X1    g368(.A1(new_n569_), .A2(KEYINPUT80), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n566_), .B(new_n570_), .Z(new_n571_));
  NOR4_X1   g370(.A1(new_n391_), .A2(new_n559_), .A3(new_n560_), .A4(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n485_), .A3(new_n313_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT100), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT100), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(KEYINPUT38), .A3(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n352_), .A2(new_n364_), .A3(new_n390_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n324_), .A2(new_n352_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n385_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n557_), .A2(new_n571_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT101), .ZN(new_n582_));
  INV_X1    g381(.A(new_n516_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n517_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G1gat), .B1(new_n585_), .B2(new_n314_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n576_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT38), .B1(new_n574_), .B2(new_n575_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(G1324gat));
  OAI21_X1  g388(.A(G8gat), .B1(new_n585_), .B2(new_n364_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT39), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n572_), .A2(new_n486_), .A3(new_n388_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(G1325gat));
  OAI21_X1  g394(.A(G15gat), .B1(new_n585_), .B2(new_n385_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT41), .Z(new_n597_));
  NAND3_X1  g396(.A1(new_n572_), .A2(new_n369_), .A3(new_n579_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(G1326gat));
  OAI21_X1  g398(.A(G22gat), .B1(new_n585_), .B2(new_n352_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT42), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n352_), .A2(G22gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT103), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n572_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(G1327gat));
  INV_X1    g404(.A(new_n571_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n517_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n557_), .A2(new_n607_), .A3(new_n516_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n580_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n609_), .A2(G29gat), .A3(new_n314_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT43), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n484_), .A2(new_n518_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n580_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n580_), .B2(new_n612_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n583_), .B(new_n582_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT44), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n482_), .A2(new_n483_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT37), .B1(new_n517_), .B2(KEYINPUT76), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT43), .B1(new_n391_), .B2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n580_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n623_), .A2(KEYINPUT44), .A3(new_n583_), .A4(new_n582_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n617_), .A2(new_n313_), .A3(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n625_), .A2(KEYINPUT104), .A3(G29gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT104), .B1(new_n625_), .B2(G29gat), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n610_), .B1(new_n626_), .B2(new_n627_), .ZN(G1328gat));
  NAND3_X1  g427(.A1(new_n617_), .A2(new_n388_), .A3(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(G36gat), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n364_), .A2(G36gat), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n609_), .A2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT45), .Z(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT46), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n630_), .A2(KEYINPUT46), .A3(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1329gat));
  NAND4_X1  g437(.A1(new_n617_), .A2(new_n624_), .A3(G43gat), .A4(new_n579_), .ZN(new_n639_));
  INV_X1    g438(.A(G43gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n609_), .B2(new_n385_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g442(.A1(new_n617_), .A2(new_n624_), .A3(G50gat), .A4(new_n351_), .ZN(new_n644_));
  INV_X1    g443(.A(G50gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n609_), .B2(new_n352_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1331gat));
  INV_X1    g446(.A(new_n557_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n606_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n580_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(new_n584_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G57gat), .B1(new_n652_), .B2(new_n314_), .ZN(new_n653_));
  NOR4_X1   g452(.A1(new_n391_), .A2(new_n648_), .A3(new_n519_), .A4(new_n606_), .ZN(new_n654_));
  INV_X1    g453(.A(G57gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n313_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(G1332gat));
  INV_X1    g456(.A(G64gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(new_n658_), .A3(new_n388_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G64gat), .B1(new_n652_), .B2(new_n364_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(KEYINPUT48), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(KEYINPUT48), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(G1333gat));
  INV_X1    g462(.A(G71gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n654_), .A2(new_n664_), .A3(new_n579_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G71gat), .B1(new_n652_), .B2(new_n385_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(KEYINPUT49), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(KEYINPUT49), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n667_), .B2(new_n668_), .ZN(G1334gat));
  INV_X1    g468(.A(G78gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n654_), .A2(new_n670_), .A3(new_n351_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G78gat), .B1(new_n652_), .B2(new_n352_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(KEYINPUT50), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(KEYINPUT50), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(G1335gat));
  NAND3_X1  g474(.A1(new_n623_), .A2(new_n583_), .A3(new_n649_), .ZN(new_n676_));
  INV_X1    g475(.A(G85gat), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n314_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n580_), .A2(new_n583_), .A3(new_n517_), .A4(new_n649_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT105), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(new_n313_), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n681_), .A2(KEYINPUT106), .A3(G85gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT106), .B1(new_n681_), .B2(G85gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n678_), .B1(new_n682_), .B2(new_n683_), .ZN(G1336gat));
  OAI21_X1  g483(.A(G92gat), .B1(new_n676_), .B2(new_n364_), .ZN(new_n685_));
  INV_X1    g484(.A(G92gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n680_), .A2(new_n686_), .A3(new_n388_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1337gat));
  OAI21_X1  g487(.A(G99gat), .B1(new_n676_), .B2(new_n385_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n579_), .A2(new_n412_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT107), .B1(new_n680_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g492(.A1(new_n680_), .A2(new_n413_), .A3(new_n351_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n623_), .A2(new_n583_), .A3(new_n351_), .A4(new_n649_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT52), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(new_n696_), .A3(G106gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n695_), .B2(G106gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT53), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT53), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n694_), .B(new_n701_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1339gat));
  XOR2_X1   g502(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT112), .B1(new_n538_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT112), .ZN(new_n706_));
  INV_X1    g505(.A(new_n704_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n544_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n541_), .B(KEYINPUT55), .C1(new_n542_), .C2(new_n543_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n528_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n529_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n705_), .A2(new_n708_), .A3(new_n709_), .A4(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(KEYINPUT56), .A3(new_n526_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT56), .B1(new_n713_), .B2(new_n526_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n547_), .B(new_n606_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n562_), .B1(new_n494_), .B2(new_n422_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n564_), .A2(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n569_), .B(new_n719_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n721_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n722_), .A2(new_n723_), .B1(new_n569_), .B2(new_n566_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n555_), .A3(new_n554_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n517_), .B1(new_n717_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT114), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT57), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT57), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n717_), .A2(new_n725_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT114), .B(new_n729_), .C1(new_n730_), .C2(new_n517_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n724_), .A2(new_n547_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n714_), .B1(new_n716_), .B2(KEYINPUT115), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n734_), .B(KEYINPUT56), .C1(new_n713_), .C2(new_n526_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n732_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT116), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT58), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT116), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n732_), .B(new_n739_), .C1(new_n733_), .C2(new_n735_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n737_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n732_), .B(KEYINPUT58), .C1(new_n733_), .C2(new_n735_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n528_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n709_), .B1(new_n746_), .B2(new_n529_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n706_), .B1(new_n544_), .B2(new_n707_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n546_), .B1(new_n749_), .B2(new_n708_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n734_), .B1(new_n750_), .B2(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n716_), .A2(KEYINPUT115), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n714_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n753_), .A2(KEYINPUT117), .A3(KEYINPUT58), .A4(new_n732_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n744_), .A2(new_n754_), .A3(new_n612_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n728_), .B(new_n731_), .C1(new_n741_), .C2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n583_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n550_), .A2(new_n556_), .A3(new_n571_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n758_), .A2(new_n516_), .A3(new_n484_), .A4(new_n518_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n759_), .A2(KEYINPUT109), .A3(KEYINPUT54), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT109), .B1(new_n759_), .B2(KEYINPUT54), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n550_), .A2(new_n556_), .A3(new_n763_), .A4(new_n571_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n620_), .A2(KEYINPUT108), .A3(new_n516_), .A4(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n519_), .B2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT110), .B1(new_n762_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n550_), .A2(new_n556_), .A3(new_n571_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT54), .B1(new_n519_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n759_), .A2(KEYINPUT109), .A3(KEYINPUT54), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n769_), .A2(new_n774_), .A3(KEYINPUT110), .A4(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n757_), .B1(new_n770_), .B2(new_n777_), .ZN(new_n778_));
  NOR4_X1   g577(.A1(new_n388_), .A2(new_n351_), .A3(new_n314_), .A4(new_n385_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(G113gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n606_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(KEYINPUT59), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n780_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n571_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n787_), .B2(new_n782_), .ZN(G1340gat));
  AOI21_X1  g587(.A(new_n648_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n789_));
  INV_X1    g588(.A(G120gat), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n648_), .A2(KEYINPUT60), .ZN(new_n791_));
  MUX2_X1   g590(.A(KEYINPUT60), .B(new_n791_), .S(new_n790_), .Z(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT118), .B1(new_n781_), .B2(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n781_), .A2(KEYINPUT118), .A3(new_n792_), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n789_), .A2(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(G1341gat));
  AOI21_X1  g594(.A(G127gat), .B1(new_n781_), .B2(new_n516_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n784_), .A2(new_n786_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n516_), .A2(G127gat), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT119), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n797_), .B2(new_n799_), .ZN(G1342gat));
  INV_X1    g599(.A(G134gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n781_), .A2(new_n801_), .A3(new_n517_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n620_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n801_), .ZN(G1343gat));
  NOR4_X1   g603(.A1(new_n388_), .A2(new_n352_), .A3(new_n314_), .A4(new_n579_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n778_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n606_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g608(.A1(new_n806_), .A2(new_n648_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT120), .B(G148gat), .Z(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(G1345gat));
  NAND3_X1  g611(.A1(new_n807_), .A2(KEYINPUT121), .A3(new_n516_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n806_), .B2(new_n583_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT61), .B(G155gat), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n813_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1346gat));
  OR3_X1    g618(.A1(new_n806_), .A2(G162gat), .A3(new_n607_), .ZN(new_n820_));
  OAI21_X1  g619(.A(G162gat), .B1(new_n806_), .B2(new_n620_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1347gat));
  INV_X1    g621(.A(KEYINPUT62), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n769_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n826_), .A2(new_n776_), .B1(new_n583_), .B2(new_n756_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n388_), .A2(new_n352_), .A3(new_n390_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n606_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n823_), .B1(new_n830_), .B2(G169gat), .ZN(new_n831_));
  AOI211_X1 g630(.A(KEYINPUT62), .B(new_n268_), .C1(new_n829_), .C2(new_n606_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n827_), .A2(KEYINPUT122), .A3(new_n828_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n834_));
  INV_X1    g633(.A(new_n828_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n778_), .B2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n571_), .A2(new_n263_), .ZN(new_n838_));
  OAI22_X1  g637(.A1(new_n831_), .A2(new_n832_), .B1(new_n837_), .B2(new_n838_), .ZN(G1348gat));
  NOR4_X1   g638(.A1(new_n827_), .A2(new_n269_), .A3(new_n648_), .A4(new_n828_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n557_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n269_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT122), .B1(new_n827_), .B2(new_n828_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n778_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n648_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT123), .B1(new_n846_), .B2(G176gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n840_), .B1(new_n843_), .B2(new_n847_), .ZN(G1349gat));
  AOI21_X1  g647(.A(G183gat), .B1(new_n829_), .B2(new_n516_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n837_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n583_), .A2(new_n265_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(G1350gat));
  OAI21_X1  g651(.A(G190gat), .B1(new_n837_), .B2(new_n620_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n517_), .A2(new_n266_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n837_), .B2(new_n854_), .ZN(G1351gat));
  AND3_X1   g654(.A1(new_n388_), .A2(new_n365_), .A3(new_n385_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n778_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n571_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n246_), .ZN(G1352gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n648_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT124), .B(G204gat), .Z(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n860_), .B2(new_n863_), .ZN(G1353gat));
  AND2_X1   g663(.A1(new_n778_), .A2(new_n856_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n866_));
  INV_X1    g665(.A(G211gat), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n865_), .B(new_n516_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n867_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT125), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n868_), .B(new_n870_), .ZN(G1354gat));
  NAND2_X1  g670(.A1(new_n612_), .A2(G218gat), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT126), .Z(new_n873_));
  NAND2_X1  g672(.A1(new_n865_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n857_), .A2(new_n607_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(G218gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT127), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT127), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n874_), .B(new_n878_), .C1(new_n875_), .C2(G218gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1355gat));
endmodule


