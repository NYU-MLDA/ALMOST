//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n862_, new_n864_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT89), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n205_));
  OR2_X1    g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(new_n207_), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n205_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT91), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(KEYINPUT91), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT22), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT90), .B1(new_n214_), .B2(G169gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT22), .B(G169gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n213_), .B(new_n215_), .C1(new_n216_), .C2(KEYINPUT90), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n213_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n212_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  AOI211_X1 g023(.A(new_n221_), .B(new_n222_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  MUX2_X1   g024(.A(new_n202_), .B(new_n204_), .S(new_n207_), .Z(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n218_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT99), .ZN(new_n230_));
  INV_X1    g029(.A(G204gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G197gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT98), .B(G197gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n232_), .B1(new_n233_), .B2(new_n231_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT21), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237_));
  OAI211_X1 g036(.A(KEYINPUT21), .B(new_n237_), .C1(new_n233_), .C2(G204gat), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n230_), .B(new_n238_), .C1(KEYINPUT21), .C2(new_n234_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n228_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT20), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n226_), .A2(new_n206_), .B1(G169gat), .B2(G176gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n216_), .A2(new_n213_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n205_), .A2(new_n208_), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n243_), .A2(new_n244_), .B1(new_n225_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n240_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n242_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G226gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT19), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G8gat), .B(G36gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT104), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G64gat), .B(G92gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT103), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n246_), .A2(new_n247_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n218_), .A2(new_n227_), .A3(new_n247_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(KEYINPUT20), .A4(new_n251_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n253_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n259_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n262_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n251_), .B1(new_n241_), .B2(new_n248_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT105), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n265_), .A2(new_n266_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(KEYINPUT105), .A3(new_n259_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G1gat), .B(G29gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT109), .ZN(new_n274_));
  XOR2_X1   g073(.A(G57gat), .B(G85gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT108), .B(KEYINPUT0), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  AND2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n279_), .B2(KEYINPUT1), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT94), .Z(new_n288_));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT95), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(new_n285_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(KEYINPUT95), .B2(new_n289_), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n284_), .B(KEYINPUT2), .Z(new_n293_));
  OAI21_X1  g092(.A(new_n281_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n288_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT93), .B(G127gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G134gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n288_), .A2(new_n299_), .A3(new_n294_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n295_), .A2(new_n308_), .A3(new_n300_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT107), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT106), .B1(new_n303_), .B2(new_n308_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT106), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n301_), .A2(new_n313_), .A3(KEYINPUT4), .A4(new_n302_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n278_), .B(new_n307_), .C1(new_n315_), .C2(new_n306_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT33), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n306_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n304_), .A2(new_n306_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n278_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n317_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n319_), .B1(new_n315_), .B2(new_n306_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n324_), .A2(KEYINPUT33), .A3(new_n278_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n272_), .B(new_n316_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT110), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n321_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT33), .B1(new_n324_), .B2(new_n278_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT110), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(new_n316_), .A4(new_n272_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n270_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT111), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n249_), .A2(new_n251_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n260_), .A2(new_n261_), .A3(KEYINPUT20), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n251_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n333_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n321_), .A2(new_n322_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n324_), .A2(new_n278_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n335_), .B(new_n339_), .C1(new_n340_), .C2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n327_), .A2(new_n332_), .A3(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT100), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n288_), .B2(new_n294_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(new_n247_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G228gat), .A2(G233gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT101), .ZN(new_n352_));
  OAI211_X1 g151(.A(G228gat), .B(G233gat), .C1(new_n348_), .C2(new_n247_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n346_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT102), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT97), .B1(new_n295_), .B2(KEYINPUT29), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n295_), .A2(KEYINPUT97), .A3(KEYINPUT29), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n359_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n359_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n363_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n351_), .A2(new_n345_), .A3(new_n353_), .ZN(new_n373_));
  OAI211_X1 g172(.A(KEYINPUT102), .B(new_n346_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n358_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n351_), .A2(new_n353_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n346_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n373_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n370_), .A2(new_n378_), .A3(new_n371_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n299_), .B(KEYINPUT92), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT31), .ZN(new_n382_));
  INV_X1    g181(.A(new_n228_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G15gat), .B(G43gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT30), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G71gat), .B(G99gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n384_), .B(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n380_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n343_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n340_), .A2(new_n341_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n391_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n380_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n391_), .A2(new_n379_), .A3(new_n375_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n272_), .A2(KEYINPUT27), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n338_), .A2(new_n259_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(KEYINPUT27), .A3(new_n267_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n393_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(KEYINPUT13), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(KEYINPUT13), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G230gat), .A2(G233gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT65), .B(G106gat), .Z(new_n411_));
  INV_X1    g210(.A(G99gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT10), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT10), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G99gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT64), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n411_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT66), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421_));
  INV_X1    g220(.A(G106gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n412_), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(G85gat), .A2(G92gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(G85gat), .A2(G92gat), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT67), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT9), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n426_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT9), .B1(new_n427_), .B2(new_n428_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n425_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT66), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n434_), .B(new_n411_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n420_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT68), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n420_), .A2(KEYINPUT68), .A3(new_n433_), .A4(new_n435_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G99gat), .A2(G106gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(KEYINPUT69), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n443_), .A2(new_n423_), .A3(new_n424_), .A4(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT70), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n427_), .A2(new_n426_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT8), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT8), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n441_), .A2(new_n442_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(KEYINPUT69), .B2(KEYINPUT7), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n423_), .A2(new_n444_), .A3(new_n424_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n450_), .B(new_n447_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n438_), .A2(new_n439_), .A3(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(G57gat), .A2(G64gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G57gat), .A2(G64gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT11), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT71), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n461_), .B(KEYINPUT11), .C1(new_n457_), .C2(new_n458_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  OR3_X1    g262(.A1(new_n457_), .A2(new_n458_), .A3(KEYINPUT11), .ZN(new_n464_));
  XOR2_X1   g263(.A(G71gat), .B(G78gat), .Z(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n460_), .A2(new_n464_), .A3(new_n465_), .A4(new_n462_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n456_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n438_), .A2(new_n439_), .A3(new_n455_), .A4(new_n469_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n410_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT72), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n454_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n450_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT73), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT73), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n449_), .A2(new_n479_), .A3(new_n454_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n438_), .A2(new_n439_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT75), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n467_), .A2(KEYINPUT74), .A3(new_n468_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT74), .B1(new_n467_), .B2(new_n468_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT12), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n481_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n482_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT12), .B1(new_n456_), .B2(new_n470_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT76), .B1(new_n472_), .B2(new_n410_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n472_), .A2(KEYINPUT76), .A3(new_n410_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n475_), .A2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G120gat), .B(G148gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G176gat), .B(G204gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n496_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT78), .B1(new_n496_), .B2(new_n502_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n475_), .A2(new_n495_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n507_), .A2(KEYINPUT78), .A3(new_n501_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n408_), .B(new_n409_), .C1(new_n506_), .C2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n501_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(KEYINPUT78), .A3(new_n503_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n510_), .A2(new_n512_), .A3(KEYINPUT79), .A4(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n509_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT80), .B(G43gat), .ZN(new_n516_));
  INV_X1    g315(.A(G50gat), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n516_), .A2(new_n517_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G29gat), .B(G36gat), .ZN(new_n520_));
  OR3_X1    g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525_));
  INV_X1    g324(.A(G1gat), .ZN(new_n526_));
  INV_X1    g325(.A(G8gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G1gat), .B(G8gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n524_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n523_), .B(KEYINPUT15), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n533_), .B2(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n523_), .B(new_n531_), .Z(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(G229gat), .A3(G233gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n536_), .B1(KEYINPUT88), .B2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(KEYINPUT88), .B2(new_n538_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(new_n219_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(G197gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n540_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n515_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n405_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n531_), .B(KEYINPUT85), .ZN(new_n548_));
  AND2_X1   g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(new_n470_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT74), .B(KEYINPUT86), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT16), .B(G183gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G211gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n553_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n553_), .A2(KEYINPUT87), .A3(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n559_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n557_), .A2(new_n558_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n551_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n533_), .A2(new_n481_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(KEYINPUT82), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT34), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(KEYINPUT35), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT81), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n571_), .B(new_n577_), .C1(new_n524_), .C2(new_n456_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n456_), .A2(new_n524_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n533_), .B2(new_n481_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n581_), .A2(new_n572_), .A3(new_n574_), .A4(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(G134gat), .ZN(new_n585_));
  INV_X1    g384(.A(G162gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n589_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n587_), .A2(new_n588_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n579_), .B(new_n582_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(KEYINPUT37), .A3(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n594_), .A2(KEYINPUT83), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(KEYINPUT83), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n590_), .A2(new_n593_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT84), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT84), .ZN(new_n600_));
  AOI211_X1 g399(.A(new_n600_), .B(KEYINPUT37), .C1(new_n590_), .C2(new_n593_), .ZN(new_n601_));
  OAI22_X1  g400(.A1(new_n595_), .A2(new_n596_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n569_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n547_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n526_), .A3(new_n395_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT38), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n547_), .A2(new_n568_), .A3(new_n597_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(new_n395_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n526_), .B2(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(new_n403_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n604_), .A2(new_n527_), .A3(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n568_), .A2(new_n597_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n405_), .A2(new_n546_), .A3(new_n610_), .A4(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n613_), .A2(new_n614_), .A3(G8gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n613_), .B2(G8gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n611_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT112), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g418(.A(G15gat), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n607_), .B2(new_n391_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT41), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n604_), .A2(new_n620_), .A3(new_n391_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1326gat));
  INV_X1    g423(.A(G22gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n607_), .B2(new_n380_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT42), .Z(new_n627_));
  NAND3_X1  g426(.A1(new_n604_), .A2(new_n625_), .A3(new_n380_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1327gat));
  AOI22_X1  g428(.A1(new_n343_), .A2(new_n392_), .B1(new_n399_), .B2(new_n403_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n515_), .A2(new_n545_), .A3(new_n568_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n597_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(G29gat), .B1(new_n633_), .B2(new_n395_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n602_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT114), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT43), .B1(new_n602_), .B2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n405_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n637_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n630_), .B2(new_n602_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT113), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n631_), .B(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(G29gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n641_), .A2(new_n643_), .A3(KEYINPUT44), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n394_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n634_), .B1(new_n647_), .B2(new_n650_), .ZN(G1328gat));
  INV_X1    g450(.A(G36gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n403_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(new_n648_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n633_), .A2(new_n652_), .A3(new_n610_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT45), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n655_), .A2(KEYINPUT115), .A3(new_n656_), .A4(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(KEYINPUT115), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n656_), .A2(KEYINPUT115), .ZN(new_n661_));
  INV_X1    g460(.A(new_n658_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n660_), .B(new_n661_), .C1(new_n654_), .C2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n659_), .A2(new_n663_), .ZN(G1329gat));
  INV_X1    g463(.A(KEYINPUT47), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n646_), .A2(G43gat), .A3(new_n391_), .A4(new_n648_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT116), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n633_), .A2(new_n391_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(G43gat), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n666_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n667_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n665_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n666_), .A2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT116), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n666_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(KEYINPUT47), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n672_), .A2(new_n676_), .ZN(G1330gat));
  AOI21_X1  g476(.A(G50gat), .B1(new_n633_), .B2(new_n380_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n380_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n649_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n517_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1331gat));
  NOR2_X1   g481(.A1(new_n515_), .A2(new_n545_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n405_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AND4_X1   g484(.A1(G57gat), .A2(new_n685_), .A3(new_n395_), .A4(new_n612_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n684_), .A2(new_n603_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT117), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT117), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n395_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(G57gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n686_), .B1(new_n690_), .B2(new_n691_), .ZN(G1332gat));
  NOR2_X1   g491(.A1(new_n403_), .A2(G64gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(new_n689_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n685_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(G64gat), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n695_), .A3(G64gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1333gat));
  NOR2_X1   g498(.A1(new_n396_), .A2(G71gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n688_), .A2(new_n689_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT49), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n685_), .A2(new_n391_), .A3(new_n612_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(G71gat), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(new_n702_), .A3(G71gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(G1334gat));
  NOR2_X1   g505(.A1(new_n679_), .A2(G78gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n688_), .A2(new_n689_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT50), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n685_), .A2(new_n380_), .A3(new_n612_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G78gat), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n709_), .A3(G78gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(G1335gat));
  NOR3_X1   g512(.A1(new_n515_), .A2(new_n545_), .A3(new_n569_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n715_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G85gat), .B1(new_n716_), .B2(new_n395_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(new_n395_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n719_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g519(.A(G92gat), .B1(new_n716_), .B2(new_n610_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n610_), .A2(G92gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n718_), .B2(new_n722_), .ZN(G1337gat));
  OAI211_X1 g522(.A(new_n716_), .B(new_n391_), .C1(new_n418_), .C2(new_n417_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n718_), .A2(new_n391_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n412_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g526(.A1(new_n716_), .A2(new_n411_), .A3(new_n380_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n718_), .A2(new_n380_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(G106gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT52), .B(new_n422_), .C1(new_n718_), .C2(new_n380_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g533(.A1(new_n509_), .A2(new_n514_), .A3(new_n544_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT54), .B1(new_n603_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n594_), .B(KEYINPUT83), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n597_), .A2(new_n598_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n600_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n597_), .A2(KEYINPUT84), .A3(new_n598_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n568_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT54), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n742_), .A2(new_n515_), .A3(new_n743_), .A4(new_n544_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n736_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n488_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n489_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n481_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n472_), .ZN(new_n750_));
  OAI211_X1 g549(.A(G230gat), .B(G233gat), .C1(new_n749_), .C2(new_n750_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n472_), .A2(KEYINPUT76), .A3(new_n410_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(new_n491_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n749_), .A2(new_n753_), .A3(KEYINPUT55), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n751_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT118), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT118), .B(new_n751_), .C1(new_n754_), .C2(new_n756_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n502_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT56), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT56), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n759_), .A2(new_n763_), .A3(new_n502_), .A4(new_n760_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n762_), .A2(new_n511_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n766_));
  MUX2_X1   g565(.A(new_n534_), .B(new_n537_), .S(new_n535_), .Z(new_n767_));
  INV_X1    g566(.A(new_n543_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n540_), .B2(new_n768_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n765_), .A2(new_n766_), .A3(KEYINPUT58), .A4(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n762_), .A2(new_n511_), .A3(new_n770_), .A4(new_n764_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT58), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n602_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT119), .B1(new_n772_), .B2(new_n773_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n771_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n762_), .A2(new_n545_), .A3(new_n511_), .A4(new_n764_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n510_), .A2(new_n512_), .A3(new_n770_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n632_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n776_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n745_), .B1(new_n784_), .B2(new_n568_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n610_), .A2(new_n394_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n785_), .A2(new_n398_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G113gat), .B1(new_n788_), .B2(new_n545_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n398_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT57), .B1(new_n779_), .B2(new_n632_), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n781_), .B(new_n597_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n569_), .B1(new_n793_), .B2(new_n776_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n790_), .B(new_n786_), .C1(new_n794_), .C2(new_n745_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT59), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n784_), .A2(new_n568_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n745_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n801_), .A2(new_n790_), .A3(new_n786_), .A4(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n544_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n789_), .B1(new_n804_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g604(.A(G120gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n515_), .B2(KEYINPUT60), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n788_), .B(new_n807_), .C1(KEYINPUT60), .C2(new_n806_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n515_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n806_), .ZN(G1341gat));
  INV_X1    g609(.A(G127gat), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n568_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n797_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n787_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n790_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n802_), .ZN(new_n816_));
  NOR4_X1   g615(.A1(new_n785_), .A2(new_n398_), .A3(new_n787_), .A4(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n812_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n811_), .B1(new_n795_), .B2(new_n568_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT121), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n812_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n822_));
  AOI21_X1  g621(.A(G127gat), .B1(new_n788_), .B2(new_n569_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n820_), .A2(new_n825_), .ZN(G1342gat));
  AOI21_X1  g625(.A(G134gat), .B1(new_n788_), .B2(new_n597_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n602_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g628(.A1(new_n785_), .A2(new_n397_), .A3(new_n787_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n545_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g631(.A(new_n515_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g634(.A1(new_n830_), .A2(new_n569_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT61), .B(G155gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1346gat));
  NAND2_X1  g637(.A1(new_n830_), .A2(new_n597_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n586_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n830_), .A2(G162gat), .A3(new_n635_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n840_), .A2(KEYINPUT122), .A3(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1347gat));
  NOR2_X1   g645(.A1(new_n403_), .A2(new_n395_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n785_), .A2(new_n398_), .A3(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT123), .A3(new_n545_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n790_), .B(new_n847_), .C1(new_n794_), .C2(new_n745_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n544_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(G169gat), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n849_), .A2(new_n545_), .A3(new_n216_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n850_), .A2(KEYINPUT62), .A3(new_n853_), .A4(G169gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(G1348gat));
  NOR2_X1   g658(.A1(new_n852_), .A2(new_n515_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n213_), .ZN(G1349gat));
  NOR2_X1   g660(.A1(new_n852_), .A2(new_n568_), .ZN(new_n862_));
  MUX2_X1   g661(.A(G183gat), .B(new_n223_), .S(new_n862_), .Z(G1350gat));
  OAI21_X1  g662(.A(G190gat), .B1(new_n852_), .B2(new_n602_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n597_), .A2(new_n224_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT124), .Z(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n852_), .B2(new_n866_), .ZN(G1351gat));
  NOR3_X1   g666(.A1(new_n785_), .A2(new_n397_), .A3(new_n848_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n545_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n833_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g671(.A1(new_n848_), .A2(new_n397_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n801_), .A2(new_n873_), .ZN(new_n874_));
  OAI22_X1  g673(.A1(new_n874_), .A2(new_n568_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT63), .B(G211gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n868_), .A2(new_n569_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1354gat));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n874_), .B2(new_n632_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n868_), .A2(KEYINPUT126), .A3(new_n597_), .ZN(new_n883_));
  INV_X1    g682(.A(G218gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n868_), .A2(G218gat), .A3(new_n635_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1355gat));
endmodule


