//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n987_, new_n988_,
    new_n989_;
  INV_X1    g000(.A(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G148gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT3), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(G141gat), .B2(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT86), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(KEYINPUT86), .A3(new_n209_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n207_), .A2(new_n212_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT85), .B1(new_n216_), .B2(KEYINPUT1), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT85), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(G155gat), .A4(G162gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(KEYINPUT1), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n219_), .A2(new_n222_), .A3(new_n217_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n202_), .A2(new_n203_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n208_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n218_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT87), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT29), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT87), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n218_), .A2(new_n230_), .A3(new_n226_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n233_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n228_), .A2(new_n229_), .A3(new_n231_), .A4(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G22gat), .B(G50gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n234_), .A2(new_n238_), .A3(new_n236_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT21), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G204gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n245_), .B2(KEYINPUT89), .ZN(new_n246_));
  INV_X1    g045(.A(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G197gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n246_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(KEYINPUT90), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT91), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G197gat), .B(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT91), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n257_), .A3(KEYINPUT21), .ZN(new_n258_));
  OAI22_X1  g057(.A1(new_n250_), .A2(new_n252_), .B1(new_n253_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT92), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI221_X1 g060(.A(KEYINPUT92), .B1(new_n253_), .B2(new_n258_), .C1(new_n250_), .C2(new_n252_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G228gat), .A2(G233gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n218_), .A2(new_n230_), .A3(new_n226_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n230_), .B1(new_n218_), .B2(new_n226_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT29), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n259_), .A3(new_n265_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G78gat), .B(G106gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT93), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT94), .Z(new_n274_));
  NAND3_X1  g073(.A1(new_n267_), .A2(new_n271_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT95), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n267_), .A2(new_n271_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n273_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n267_), .A2(new_n271_), .A3(KEYINPUT95), .A4(new_n274_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n242_), .A2(new_n277_), .A3(new_n279_), .A4(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n275_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n274_), .B1(new_n267_), .B2(new_n271_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n241_), .B(new_n240_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G183gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT79), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G183gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT80), .ZN(new_n290_));
  OAI211_X1 g089(.A(KEYINPUT25), .B(new_n287_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n291_));
  OR3_X1    g090(.A1(new_n290_), .A2(new_n286_), .A3(KEYINPUT25), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G190gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT81), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(G176gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n294_), .A2(KEYINPUT81), .B1(KEYINPUT24), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT23), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(G183gat), .A3(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(KEYINPUT24), .B2(new_n298_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT82), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n309_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n295_), .A2(new_n302_), .A3(new_n310_), .A4(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n287_), .A2(new_n289_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n307_), .B1(new_n313_), .B2(G190gat), .ZN(new_n314_));
  OR2_X1    g113(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n297_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n299_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT84), .B(G113gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G120gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(G127gat), .B(G134gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n323_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n322_), .B(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n312_), .A2(new_n327_), .A3(new_n319_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G71gat), .B(G99gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT31), .ZN(new_n333_));
  XOR2_X1   g132(.A(G15gat), .B(G43gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G227gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n325_), .A2(new_n328_), .A3(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n331_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n331_), .B2(new_n339_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n285_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n340_), .A2(new_n341_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n327_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT99), .B1(new_n347_), .B2(KEYINPUT4), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n324_), .A2(new_n226_), .A3(new_n218_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n349_), .A3(KEYINPUT4), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n228_), .A2(new_n231_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT99), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .A4(new_n327_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n348_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT101), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT0), .B(G57gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G85gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(G1gat), .B(G29gat), .Z(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n358_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT102), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n359_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT101), .B1(new_n371_), .B2(new_n366_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT102), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n373_), .A3(new_n366_), .ZN(new_n374_));
  AND4_X1   g173(.A1(new_n368_), .A2(new_n370_), .A3(new_n372_), .A4(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT18), .B(G64gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G92gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT19), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n261_), .A2(new_n262_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n300_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT25), .B(G183gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n293_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n386_), .A2(new_n388_), .A3(new_n307_), .A4(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n286_), .A2(new_n391_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n307_), .A2(new_n392_), .B1(new_n317_), .B2(new_n297_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n299_), .B(KEYINPUT97), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n384_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n320_), .B2(new_n259_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n383_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n253_), .A2(new_n258_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n246_), .A2(new_n256_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n246_), .A2(new_n256_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n252_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n312_), .A2(new_n404_), .A3(new_n319_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT98), .B1(new_n393_), .B2(new_n394_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n307_), .A2(new_n392_), .ZN(new_n407_));
  AND4_X1   g206(.A1(KEYINPUT98), .A2(new_n407_), .A3(new_n318_), .A4(new_n394_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n390_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n259_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n405_), .A2(new_n411_), .A3(KEYINPUT20), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n412_), .A2(new_n382_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n380_), .B1(new_n399_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n382_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n409_), .A2(new_n410_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n382_), .B1(new_n416_), .B2(new_n404_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n398_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n418_), .A3(new_n379_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n414_), .A2(KEYINPUT27), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT27), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n415_), .A2(new_n418_), .A3(new_n379_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n379_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT103), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT103), .B(new_n421_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n420_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n346_), .A2(new_n375_), .A3(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n368_), .A2(new_n370_), .A3(new_n372_), .A4(new_n374_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n379_), .A2(KEYINPUT32), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n415_), .A2(new_n418_), .A3(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n432_), .B(KEYINPUT100), .Z(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT32), .B(new_n379_), .C1(new_n399_), .C2(new_n413_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n422_), .A2(new_n423_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n347_), .A2(new_n349_), .A3(new_n357_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n366_), .B(new_n437_), .C1(new_n355_), .C2(new_n357_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n361_), .A2(new_n367_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n440_), .A2(KEYINPUT33), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(KEYINPUT33), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n344_), .B1(new_n435_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n285_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n429_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G113gat), .B(G141gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(new_n296_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(G197gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G229gat), .A2(G233gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G1gat), .A2(G8gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT14), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT73), .ZN(new_n455_));
  OR2_X1    g254(.A1(G15gat), .A2(G22gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G15gat), .A2(G22gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT73), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n459_), .A3(KEYINPUT14), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n455_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n453_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G1gat), .A2(G8gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT74), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(G1gat), .ZN(new_n465_));
  INV_X1    g264(.A(G8gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT74), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n453_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n461_), .A2(new_n470_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(KEYINPUT73), .A2(new_n454_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n472_), .A2(new_n464_), .A3(new_n469_), .A4(new_n460_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G29gat), .A2(G36gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(G29gat), .A2(G36gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(G43gat), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G29gat), .ZN(new_n479_));
  INV_X1    g278(.A(G36gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G43gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n475_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n478_), .A2(new_n483_), .A3(G50gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(G50gat), .B1(new_n478_), .B2(new_n483_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n474_), .A2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n471_), .B(new_n473_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n487_), .A2(KEYINPUT77), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT77), .B1(new_n487_), .B2(new_n488_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n452_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n478_), .A2(new_n483_), .ZN(new_n494_));
  INV_X1    g293(.A(G50gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n478_), .A2(new_n483_), .A3(G50gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(KEYINPUT15), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n451_), .B(new_n487_), .C1(new_n500_), .C2(new_n474_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n491_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT78), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n450_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AOI211_X1 g303(.A(KEYINPUT78), .B(new_n449_), .C1(new_n491_), .C2(new_n501_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT13), .ZN(new_n507_));
  XOR2_X1   g306(.A(G120gat), .B(G148gat), .Z(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G176gat), .B(G204gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G99gat), .ZN(new_n517_));
  INV_X1    g316(.A(G106gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT65), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT7), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n521_), .A2(new_n517_), .A3(new_n518_), .A4(KEYINPUT65), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n516_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G85gat), .B(G92gat), .Z(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT66), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n523_), .A2(new_n524_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT10), .B(G99gat), .Z(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n518_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n524_), .A2(KEYINPUT9), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(G85gat), .A3(G92gat), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .A4(new_n516_), .ZN(new_n537_));
  INV_X1    g336(.A(G57gat), .ZN(new_n538_));
  INV_X1    g337(.A(G64gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT11), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G57gat), .A2(G64gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544_));
  OR2_X1    g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT67), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n540_), .A2(new_n542_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(new_n541_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT67), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n543_), .A2(new_n550_), .A3(new_n544_), .A4(new_n545_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n549_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n531_), .B(new_n537_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n523_), .A2(new_n524_), .A3(new_n529_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n529_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n537_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n554_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n552_), .A3(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(new_n560_), .A3(KEYINPUT12), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n553_), .A2(new_n554_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n558_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT64), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n555_), .B2(new_n560_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n513_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n567_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n573_), .A2(new_n570_), .A3(new_n512_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n507_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n569_), .A2(new_n571_), .A3(new_n513_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n512_), .B1(new_n573_), .B2(new_n570_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(KEYINPUT13), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT16), .B(G183gat), .ZN(new_n580_));
  INV_X1    g379(.A(G211gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G127gat), .B(G155gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n580_), .B(G211gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(new_n583_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT17), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n583_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n582_), .A2(new_n584_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(G231gat), .ZN(new_n594_));
  INV_X1    g393(.A(G233gat), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n474_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n471_), .A2(new_n473_), .A3(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n559_), .A2(new_n597_), .A3(new_n552_), .A4(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n598_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n602_));
  OAI22_X1  g401(.A1(new_n601_), .A2(new_n602_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n593_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n588_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n600_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT75), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n603_), .A2(new_n600_), .A3(new_n605_), .A4(KEYINPUT75), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n604_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(KEYINPUT76), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT76), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n612_), .B(new_n604_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR4_X1   g414(.A1(new_n446_), .A2(new_n506_), .A3(new_n579_), .A4(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n558_), .A2(new_n499_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT34), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT35), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n486_), .B(new_n537_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n617_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n620_), .A2(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(G134gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(G162gat), .ZN(new_n629_));
  INV_X1    g428(.A(G134gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n627_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(G162gat), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n629_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n625_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n617_), .A2(new_n637_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n626_), .A2(new_n636_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT69), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT69), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n626_), .A2(new_n641_), .A3(new_n638_), .A4(new_n636_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n634_), .B1(new_n629_), .B2(new_n633_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(KEYINPUT70), .A3(new_n635_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT70), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n647_), .B1(new_n636_), .B2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n624_), .A2(new_n625_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n638_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT71), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n649_), .B1(new_n626_), .B2(new_n638_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT71), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n643_), .A2(new_n654_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT37), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT72), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n626_), .A2(KEYINPUT72), .A3(new_n638_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n650_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT37), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n643_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n659_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n616_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n465_), .A3(new_n430_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT38), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n663_), .A2(new_n643_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n616_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G1gat), .B1(new_n672_), .B2(new_n375_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n673_), .ZN(G1324gat));
  INV_X1    g473(.A(new_n428_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n667_), .A2(new_n466_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT39), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n671_), .A2(new_n675_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(G8gat), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT39), .B(new_n466_), .C1(new_n671_), .C2(new_n675_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1325gat));
  INV_X1    g482(.A(new_n667_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n684_), .A2(G15gat), .A3(new_n342_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G15gat), .B1(new_n672_), .B2(new_n342_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n686_), .A2(new_n687_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(G1326gat));
  OR3_X1    g489(.A1(new_n684_), .A2(G22gat), .A3(new_n445_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G22gat), .B1(new_n672_), .B2(new_n445_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(KEYINPUT42), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(KEYINPUT42), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(G1327gat));
  NOR3_X1   g494(.A1(new_n579_), .A2(new_n506_), .A3(new_n614_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n435_), .A2(new_n443_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n445_), .A3(new_n342_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n429_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n666_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n697_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT43), .B(new_n666_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n696_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n696_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n446_), .B2(new_n666_), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n285_), .B(new_n344_), .C1(new_n435_), .C2(new_n443_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n697_), .B(new_n702_), .C1(new_n710_), .C2(new_n429_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n707_), .A2(new_n713_), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n714_), .A2(KEYINPUT104), .A3(new_n375_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT104), .B1(new_n714_), .B2(new_n375_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(G29gat), .A3(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n446_), .A2(new_n670_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n696_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n670_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n701_), .A2(new_n721_), .A3(new_n696_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT105), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n720_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n479_), .A3(new_n430_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n717_), .A2(new_n725_), .ZN(G1328gat));
  NAND4_X1  g525(.A1(new_n720_), .A2(new_n723_), .A3(new_n480_), .A4(new_n675_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT45), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n714_), .A2(new_n428_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n480_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n728_), .B(KEYINPUT46), .C1(new_n729_), .C2(new_n480_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1329gat));
  NOR2_X1   g533(.A1(new_n342_), .A2(new_n482_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n707_), .A2(new_n713_), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n720_), .A2(new_n723_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n482_), .B1(new_n738_), .B2(new_n342_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n736_), .A2(new_n737_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n736_), .B2(new_n739_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n740_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n712_), .A2(KEYINPUT44), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n706_), .B(new_n708_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n735_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n744_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G43gat), .B1(new_n724_), .B2(new_n344_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT106), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n736_), .A2(new_n737_), .A3(new_n739_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT47), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n743_), .A2(new_n751_), .ZN(G1330gat));
  OAI21_X1  g551(.A(G50gat), .B1(new_n714_), .B2(new_n445_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n724_), .A2(new_n495_), .A3(new_n285_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1331gat));
  INV_X1    g554(.A(new_n506_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n579_), .ZN(new_n757_));
  NOR4_X1   g556(.A1(new_n446_), .A2(new_n756_), .A3(new_n757_), .A4(new_n615_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n670_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(new_n538_), .A3(new_n375_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n666_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n430_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n538_), .B2(new_n763_), .ZN(G1332gat));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n539_), .A3(new_n675_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G64gat), .B1(new_n759_), .B2(new_n428_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n765_), .B1(new_n767_), .B2(new_n768_), .ZN(G1333gat));
  OR3_X1    g568(.A1(new_n761_), .A2(G71gat), .A3(new_n342_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G71gat), .B1(new_n759_), .B2(new_n342_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT49), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT49), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n772_), .B2(new_n773_), .ZN(G1334gat));
  OR3_X1    g573(.A1(new_n761_), .A2(G78gat), .A3(new_n445_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G78gat), .B1(new_n759_), .B2(new_n445_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n776_), .A2(KEYINPUT107), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(KEYINPUT107), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(KEYINPUT50), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT50), .B1(new_n777_), .B2(new_n778_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n775_), .B1(new_n779_), .B2(new_n780_), .ZN(G1335gat));
  NOR3_X1   g580(.A1(new_n757_), .A2(new_n756_), .A3(new_n614_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n718_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n430_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n709_), .A2(new_n711_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n782_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n430_), .A2(G85gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n784_), .B1(new_n788_), .B2(new_n789_), .ZN(G1336gat));
  AOI21_X1  g589(.A(G92gat), .B1(new_n783_), .B2(new_n675_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n675_), .A2(G92gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n788_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT109), .ZN(G1337gat));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n783_), .A2(new_n532_), .A3(new_n344_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n788_), .A2(new_n344_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n795_), .B(new_n796_), .C1(new_n797_), .C2(new_n517_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n517_), .B1(new_n788_), .B2(new_n344_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n796_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT51), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n783_), .A2(new_n518_), .A3(new_n285_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT110), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n785_), .A2(new_n285_), .A3(new_n782_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(G106gat), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(KEYINPUT111), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(KEYINPUT111), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n807_), .A2(KEYINPUT111), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n805_), .A2(G106gat), .A3(new_n809_), .A4(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n804_), .A2(new_n808_), .A3(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n804_), .A2(new_n813_), .A3(new_n808_), .A4(new_n811_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1339gat));
  AND3_X1   g616(.A1(new_n614_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n666_), .A2(new_n818_), .A3(new_n819_), .A4(new_n506_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n665_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n640_), .A2(new_n642_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n664_), .B1(new_n824_), .B2(new_n654_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n506_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n818_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT54), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n756_), .B1(new_n659_), .B2(new_n665_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(KEYINPUT113), .A3(new_n819_), .A4(new_n818_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n822_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n491_), .A2(new_n501_), .A3(new_n449_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n489_), .A2(new_n490_), .A3(new_n452_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n487_), .B1(new_n500_), .B2(new_n474_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n452_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n836_), .B2(new_n449_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n577_), .B2(new_n576_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n561_), .A2(new_n567_), .A3(new_n564_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT115), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n561_), .A2(new_n842_), .A3(new_n567_), .A4(new_n564_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n573_), .A2(KEYINPUT55), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n846_), .B(new_n567_), .C1(new_n561_), .C2(new_n564_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n844_), .A2(new_n845_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n839_), .B1(new_n848_), .B2(new_n513_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n569_), .A2(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n573_), .A2(KEYINPUT55), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(new_n841_), .A4(new_n843_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT56), .A3(new_n512_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n506_), .B2(new_n574_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n576_), .B(KEYINPUT114), .C1(new_n505_), .C2(new_n504_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n838_), .B1(new_n854_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n832_), .B1(new_n859_), .B2(new_n721_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(new_n857_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n849_), .B2(new_n853_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT57), .B(new_n670_), .C1(new_n862_), .C2(new_n838_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n837_), .A2(new_n574_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n852_), .A2(KEYINPUT56), .A3(new_n512_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT56), .B1(new_n852_), .B2(new_n512_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n854_), .A2(KEYINPUT58), .A3(new_n864_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n702_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n860_), .A2(new_n863_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n831_), .B1(new_n872_), .B2(new_n615_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n675_), .A2(new_n375_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n345_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n873_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877_), .B2(new_n756_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(KEYINPUT59), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n860_), .A2(new_n881_), .A3(new_n871_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n863_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n860_), .B2(new_n871_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n615_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n831_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n876_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT116), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n888_), .A2(KEYINPUT116), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n880_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n506_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n878_), .B1(new_n894_), .B2(G113gat), .ZN(G1340gat));
  XOR2_X1   g694(.A(KEYINPUT118), .B(G120gat), .Z(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n893_), .B2(new_n757_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n896_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n757_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT119), .B1(new_n898_), .B2(KEYINPUT60), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n877_), .B(new_n901_), .C1(new_n902_), .C2(new_n899_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n897_), .A2(new_n903_), .ZN(G1341gat));
  AOI21_X1  g703(.A(G127gat), .B1(new_n877_), .B2(new_n614_), .ZN(new_n905_));
  INV_X1    g704(.A(G127gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n893_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n907_), .B2(new_n614_), .ZN(G1342gat));
  AOI21_X1  g707(.A(G134gat), .B1(new_n877_), .B2(new_n721_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n893_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n666_), .A2(new_n630_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT120), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n909_), .B1(new_n910_), .B2(new_n912_), .ZN(G1343gat));
  NOR2_X1   g712(.A1(new_n873_), .A2(new_n343_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n874_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n506_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n202_), .ZN(G1344gat));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n757_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n203_), .ZN(G1345gat));
  NOR2_X1   g718(.A1(new_n915_), .A2(new_n615_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT61), .B(G155gat), .Z(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1346gat));
  NOR3_X1   g721(.A1(new_n915_), .A2(new_n632_), .A3(new_n666_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n914_), .A2(new_n721_), .A3(new_n874_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n632_), .B2(new_n924_), .ZN(G1347gat));
  AOI21_X1  g724(.A(new_n345_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n428_), .A2(new_n430_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n756_), .A2(new_n317_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n926_), .A2(new_n756_), .A3(new_n928_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n934_), .A2(new_n935_), .A3(G169gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n934_), .B2(G169gat), .ZN(new_n937_));
  OAI22_X1  g736(.A1(new_n932_), .A2(new_n933_), .B1(new_n936_), .B2(new_n937_), .ZN(G1348gat));
  NOR2_X1   g737(.A1(new_n873_), .A2(new_n285_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n939_), .A2(G176gat), .A3(new_n579_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n928_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n940_), .A2(new_n342_), .A3(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n579_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n297_), .ZN(G1349gat));
  NOR3_X1   g743(.A1(new_n941_), .A2(new_n342_), .A3(new_n615_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n313_), .B1(new_n939_), .B2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n926_), .A2(new_n928_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(KEYINPUT121), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n387_), .B1(new_n948_), .B2(new_n929_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n946_), .B1(new_n949_), .B2(new_n614_), .ZN(G1350gat));
  AOI21_X1  g749(.A(new_n666_), .B1(new_n948_), .B2(new_n929_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n721_), .A2(new_n293_), .ZN(new_n952_));
  OAI22_X1  g751(.A1(new_n951_), .A2(new_n391_), .B1(new_n932_), .B2(new_n952_), .ZN(G1351gat));
  NAND2_X1  g752(.A1(new_n872_), .A2(new_n615_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n886_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n343_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n928_), .A2(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(KEYINPUT122), .B1(new_n955_), .B2(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n873_), .A2(new_n960_), .A3(new_n957_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n959_), .A2(new_n961_), .ZN(new_n962_));
  OAI22_X1  g761(.A1(new_n962_), .A2(new_n506_), .B1(KEYINPUT123), .B2(new_n244_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n244_), .A2(KEYINPUT123), .ZN(new_n964_));
  XOR2_X1   g763(.A(new_n963_), .B(new_n964_), .Z(G1352gat));
  NOR2_X1   g764(.A1(new_n962_), .A2(new_n757_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n967_));
  AND2_X1   g766(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n966_), .B1(new_n967_), .B2(new_n968_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n969_), .B1(new_n966_), .B2(new_n967_), .ZN(G1353gat));
  OAI21_X1  g769(.A(new_n614_), .B1(new_n959_), .B2(new_n961_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n972_));
  AOI21_X1  g771(.A(KEYINPUT125), .B1(new_n971_), .B2(new_n972_), .ZN(new_n973_));
  XOR2_X1   g772(.A(KEYINPUT63), .B(G211gat), .Z(new_n974_));
  OAI211_X1 g773(.A(new_n614_), .B(new_n974_), .C1(new_n959_), .C2(new_n961_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(KEYINPUT126), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n955_), .A2(KEYINPUT122), .A3(new_n958_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n960_), .B1(new_n873_), .B2(new_n957_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n977_), .A2(new_n978_), .ZN(new_n979_));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n980_));
  NAND4_X1  g779(.A1(new_n979_), .A2(new_n980_), .A3(new_n614_), .A4(new_n974_), .ZN(new_n981_));
  AND3_X1   g780(.A1(new_n973_), .A2(new_n976_), .A3(new_n981_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n971_), .A2(new_n972_), .ZN(new_n983_));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n984_));
  AOI22_X1  g783(.A1(new_n976_), .A2(new_n981_), .B1(new_n983_), .B2(new_n984_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n982_), .A2(new_n985_), .ZN(G1354gat));
  AOI21_X1  g785(.A(G218gat), .B1(new_n979_), .B2(new_n721_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n702_), .A2(G218gat), .ZN(new_n988_));
  XOR2_X1   g787(.A(new_n988_), .B(KEYINPUT127), .Z(new_n989_));
  AOI21_X1  g788(.A(new_n987_), .B1(new_n979_), .B2(new_n989_), .ZN(G1355gat));
endmodule


